magic
tech sky130A
magscale 1 2
timestamp 1623926019
<< obsli1 >>
rect 1380 1071 118588 98481
<< obsm1 >>
rect 474 1040 119494 98592
<< metal2 >>
rect 478 99200 534 100000
rect 1398 99200 1454 100000
rect 2410 99200 2466 100000
rect 3422 99200 3478 100000
rect 4434 99200 4490 100000
rect 5446 99200 5502 100000
rect 6458 99200 6514 100000
rect 7470 99200 7526 100000
rect 8390 99200 8446 100000
rect 9402 99200 9458 100000
rect 10414 99200 10470 100000
rect 11426 99200 11482 100000
rect 12438 99200 12494 100000
rect 13450 99200 13506 100000
rect 14462 99200 14518 100000
rect 15474 99200 15530 100000
rect 16394 99200 16450 100000
rect 17406 99200 17462 100000
rect 18418 99200 18474 100000
rect 19430 99200 19486 100000
rect 20442 99200 20498 100000
rect 21454 99200 21510 100000
rect 22466 99200 22522 100000
rect 23386 99200 23442 100000
rect 24398 99200 24454 100000
rect 25410 99200 25466 100000
rect 26422 99200 26478 100000
rect 27434 99200 27490 100000
rect 28446 99200 28502 100000
rect 29458 99200 29514 100000
rect 30470 99200 30526 100000
rect 31390 99200 31446 100000
rect 32402 99200 32458 100000
rect 33414 99200 33470 100000
rect 34426 99200 34482 100000
rect 35438 99200 35494 100000
rect 36450 99200 36506 100000
rect 37462 99200 37518 100000
rect 38382 99200 38438 100000
rect 39394 99200 39450 100000
rect 40406 99200 40462 100000
rect 41418 99200 41474 100000
rect 42430 99200 42486 100000
rect 43442 99200 43498 100000
rect 44454 99200 44510 100000
rect 45466 99200 45522 100000
rect 46386 99200 46442 100000
rect 47398 99200 47454 100000
rect 48410 99200 48466 100000
rect 49422 99200 49478 100000
rect 50434 99200 50490 100000
rect 51446 99200 51502 100000
rect 52458 99200 52514 100000
rect 53378 99200 53434 100000
rect 54390 99200 54446 100000
rect 55402 99200 55458 100000
rect 56414 99200 56470 100000
rect 57426 99200 57482 100000
rect 58438 99200 58494 100000
rect 59450 99200 59506 100000
rect 60462 99200 60518 100000
rect 61382 99200 61438 100000
rect 62394 99200 62450 100000
rect 63406 99200 63462 100000
rect 64418 99200 64474 100000
rect 65430 99200 65486 100000
rect 66442 99200 66498 100000
rect 67454 99200 67510 100000
rect 68374 99200 68430 100000
rect 69386 99200 69442 100000
rect 70398 99200 70454 100000
rect 71410 99200 71466 100000
rect 72422 99200 72478 100000
rect 73434 99200 73490 100000
rect 74446 99200 74502 100000
rect 75458 99200 75514 100000
rect 76378 99200 76434 100000
rect 77390 99200 77446 100000
rect 78402 99200 78458 100000
rect 79414 99200 79470 100000
rect 80426 99200 80482 100000
rect 81438 99200 81494 100000
rect 82450 99200 82506 100000
rect 83370 99200 83426 100000
rect 84382 99200 84438 100000
rect 85394 99200 85450 100000
rect 86406 99200 86462 100000
rect 87418 99200 87474 100000
rect 88430 99200 88486 100000
rect 89442 99200 89498 100000
rect 90454 99200 90510 100000
rect 91374 99200 91430 100000
rect 92386 99200 92442 100000
rect 93398 99200 93454 100000
rect 94410 99200 94466 100000
rect 95422 99200 95478 100000
rect 96434 99200 96490 100000
rect 97446 99200 97502 100000
rect 98366 99200 98422 100000
rect 99378 99200 99434 100000
rect 100390 99200 100446 100000
rect 101402 99200 101458 100000
rect 102414 99200 102470 100000
rect 103426 99200 103482 100000
rect 104438 99200 104494 100000
rect 105450 99200 105506 100000
rect 106370 99200 106426 100000
rect 107382 99200 107438 100000
rect 108394 99200 108450 100000
rect 109406 99200 109462 100000
rect 110418 99200 110474 100000
rect 111430 99200 111486 100000
rect 112442 99200 112498 100000
rect 113362 99200 113418 100000
rect 114374 99200 114430 100000
rect 115386 99200 115442 100000
rect 116398 99200 116454 100000
rect 117410 99200 117466 100000
rect 118422 99200 118478 100000
rect 119434 99200 119490 100000
<< obsm2 >>
rect 590 99144 1342 99200
rect 1510 99144 2354 99200
rect 2522 99144 3366 99200
rect 3534 99144 4378 99200
rect 4546 99144 5390 99200
rect 5558 99144 6402 99200
rect 6570 99144 7414 99200
rect 7582 99144 8334 99200
rect 8502 99144 9346 99200
rect 9514 99144 10358 99200
rect 10526 99144 11370 99200
rect 11538 99144 12382 99200
rect 12550 99144 13394 99200
rect 13562 99144 14406 99200
rect 14574 99144 15418 99200
rect 15586 99144 16338 99200
rect 16506 99144 17350 99200
rect 17518 99144 18362 99200
rect 18530 99144 19374 99200
rect 19542 99144 20386 99200
rect 20554 99144 21398 99200
rect 21566 99144 22410 99200
rect 22578 99144 23330 99200
rect 23498 99144 24342 99200
rect 24510 99144 25354 99200
rect 25522 99144 26366 99200
rect 26534 99144 27378 99200
rect 27546 99144 28390 99200
rect 28558 99144 29402 99200
rect 29570 99144 30414 99200
rect 30582 99144 31334 99200
rect 31502 99144 32346 99200
rect 32514 99144 33358 99200
rect 33526 99144 34370 99200
rect 34538 99144 35382 99200
rect 35550 99144 36394 99200
rect 36562 99144 37406 99200
rect 37574 99144 38326 99200
rect 38494 99144 39338 99200
rect 39506 99144 40350 99200
rect 40518 99144 41362 99200
rect 41530 99144 42374 99200
rect 42542 99144 43386 99200
rect 43554 99144 44398 99200
rect 44566 99144 45410 99200
rect 45578 99144 46330 99200
rect 46498 99144 47342 99200
rect 47510 99144 48354 99200
rect 48522 99144 49366 99200
rect 49534 99144 50378 99200
rect 50546 99144 51390 99200
rect 51558 99144 52402 99200
rect 52570 99144 53322 99200
rect 53490 99144 54334 99200
rect 54502 99144 55346 99200
rect 55514 99144 56358 99200
rect 56526 99144 57370 99200
rect 57538 99144 58382 99200
rect 58550 99144 59394 99200
rect 59562 99144 60406 99200
rect 60574 99144 61326 99200
rect 61494 99144 62338 99200
rect 62506 99144 63350 99200
rect 63518 99144 64362 99200
rect 64530 99144 65374 99200
rect 65542 99144 66386 99200
rect 66554 99144 67398 99200
rect 67566 99144 68318 99200
rect 68486 99144 69330 99200
rect 69498 99144 70342 99200
rect 70510 99144 71354 99200
rect 71522 99144 72366 99200
rect 72534 99144 73378 99200
rect 73546 99144 74390 99200
rect 74558 99144 75402 99200
rect 75570 99144 76322 99200
rect 76490 99144 77334 99200
rect 77502 99144 78346 99200
rect 78514 99144 79358 99200
rect 79526 99144 80370 99200
rect 80538 99144 81382 99200
rect 81550 99144 82394 99200
rect 82562 99144 83314 99200
rect 83482 99144 84326 99200
rect 84494 99144 85338 99200
rect 85506 99144 86350 99200
rect 86518 99144 87362 99200
rect 87530 99144 88374 99200
rect 88542 99144 89386 99200
rect 89554 99144 90398 99200
rect 90566 99144 91318 99200
rect 91486 99144 92330 99200
rect 92498 99144 93342 99200
rect 93510 99144 94354 99200
rect 94522 99144 95366 99200
rect 95534 99144 96378 99200
rect 96546 99144 97390 99200
rect 97558 99144 98310 99200
rect 98478 99144 99322 99200
rect 99490 99144 100334 99200
rect 100502 99144 101346 99200
rect 101514 99144 102358 99200
rect 102526 99144 103370 99200
rect 103538 99144 104382 99200
rect 104550 99144 105394 99200
rect 105562 99144 106314 99200
rect 106482 99144 107326 99200
rect 107494 99144 108338 99200
rect 108506 99144 109350 99200
rect 109518 99144 110362 99200
rect 110530 99144 111374 99200
rect 111542 99144 112386 99200
rect 112554 99144 113306 99200
rect 113474 99144 114318 99200
rect 114486 99144 115330 99200
rect 115498 99144 116342 99200
rect 116510 99144 117354 99200
rect 117522 99144 118366 99200
rect 118534 99144 119378 99200
rect 480 1040 119488 99144
<< metal3 >>
rect 119200 87320 120000 87440
rect 119200 62296 120000 62416
rect 119200 37272 120000 37392
rect 119200 12384 120000 12504
<< obsm3 >>
rect 4484 87520 119200 98497
rect 4484 87240 119120 87520
rect 4484 62496 119200 87240
rect 4484 62216 119120 62496
rect 4484 37472 119200 62216
rect 4484 37192 119120 37472
rect 4484 12584 119200 37192
rect 4484 12304 119120 12584
rect 4484 1055 119200 12304
<< metal4 >>
rect 4484 1040 4804 98512
rect 19844 1040 20164 98512
rect 35204 1040 35524 98512
rect 50564 1040 50884 98512
rect 65924 1040 66244 98512
rect 81284 1040 81604 98512
rect 96644 1040 96964 98512
rect 112004 1040 112324 98512
<< obsm4 >>
rect 48083 95643 48149 95981
<< metal5 >>
rect 1380 96118 118588 96438
rect 1380 80800 118588 81120
rect 1380 65482 118588 65802
rect 1380 50164 118588 50484
rect 1380 34846 118588 35166
rect 1380 19528 118588 19848
rect 1380 4210 118588 4530
<< labels >>
rlabel metal3 s 119200 62296 120000 62416 6 events_o[0]
port 1 nsew signal output
rlabel metal3 s 119200 87320 120000 87440 6 events_o[1]
port 2 nsew signal output
rlabel metal3 s 119200 12384 120000 12504 6 mclk
port 3 nsew signal input
rlabel metal3 s 119200 37272 120000 37392 6 rst_n
port 4 nsew signal input
rlabel metal2 s 2410 99200 2466 100000 6 spi_clk
port 5 nsew signal output
rlabel metal2 s 3422 99200 3478 100000 6 spi_csn0
port 6 nsew signal output
rlabel metal2 s 4434 99200 4490 100000 6 spi_csn1
port 7 nsew signal output
rlabel metal2 s 5446 99200 5502 100000 6 spi_csn2
port 8 nsew signal output
rlabel metal2 s 6458 99200 6514 100000 6 spi_csn3
port 9 nsew signal output
rlabel metal2 s 7470 99200 7526 100000 6 spi_en_tx
port 10 nsew signal output
rlabel metal2 s 478 99200 534 100000 6 spi_mode[0]
port 11 nsew signal output
rlabel metal2 s 1398 99200 1454 100000 6 spi_mode[1]
port 12 nsew signal output
rlabel metal2 s 8390 99200 8446 100000 6 spi_sdi0
port 13 nsew signal input
rlabel metal2 s 9402 99200 9458 100000 6 spi_sdi1
port 14 nsew signal input
rlabel metal2 s 10414 99200 10470 100000 6 spi_sdi2
port 15 nsew signal input
rlabel metal2 s 11426 99200 11482 100000 6 spi_sdi3
port 16 nsew signal input
rlabel metal2 s 12438 99200 12494 100000 6 spi_sdo0
port 17 nsew signal output
rlabel metal2 s 13450 99200 13506 100000 6 spi_sdo1
port 18 nsew signal output
rlabel metal2 s 14462 99200 14518 100000 6 spi_sdo2
port 19 nsew signal output
rlabel metal2 s 15474 99200 15530 100000 6 spi_sdo3
port 20 nsew signal output
rlabel metal2 s 118422 99200 118478 100000 6 wbd_ack_o
port 21 nsew signal output
rlabel metal2 s 18418 99200 18474 100000 6 wbd_adr_i[0]
port 22 nsew signal input
rlabel metal2 s 28446 99200 28502 100000 6 wbd_adr_i[10]
port 23 nsew signal input
rlabel metal2 s 29458 99200 29514 100000 6 wbd_adr_i[11]
port 24 nsew signal input
rlabel metal2 s 30470 99200 30526 100000 6 wbd_adr_i[12]
port 25 nsew signal input
rlabel metal2 s 31390 99200 31446 100000 6 wbd_adr_i[13]
port 26 nsew signal input
rlabel metal2 s 32402 99200 32458 100000 6 wbd_adr_i[14]
port 27 nsew signal input
rlabel metal2 s 33414 99200 33470 100000 6 wbd_adr_i[15]
port 28 nsew signal input
rlabel metal2 s 34426 99200 34482 100000 6 wbd_adr_i[16]
port 29 nsew signal input
rlabel metal2 s 35438 99200 35494 100000 6 wbd_adr_i[17]
port 30 nsew signal input
rlabel metal2 s 36450 99200 36506 100000 6 wbd_adr_i[18]
port 31 nsew signal input
rlabel metal2 s 37462 99200 37518 100000 6 wbd_adr_i[19]
port 32 nsew signal input
rlabel metal2 s 19430 99200 19486 100000 6 wbd_adr_i[1]
port 33 nsew signal input
rlabel metal2 s 38382 99200 38438 100000 6 wbd_adr_i[20]
port 34 nsew signal input
rlabel metal2 s 39394 99200 39450 100000 6 wbd_adr_i[21]
port 35 nsew signal input
rlabel metal2 s 40406 99200 40462 100000 6 wbd_adr_i[22]
port 36 nsew signal input
rlabel metal2 s 41418 99200 41474 100000 6 wbd_adr_i[23]
port 37 nsew signal input
rlabel metal2 s 42430 99200 42486 100000 6 wbd_adr_i[24]
port 38 nsew signal input
rlabel metal2 s 43442 99200 43498 100000 6 wbd_adr_i[25]
port 39 nsew signal input
rlabel metal2 s 44454 99200 44510 100000 6 wbd_adr_i[26]
port 40 nsew signal input
rlabel metal2 s 45466 99200 45522 100000 6 wbd_adr_i[27]
port 41 nsew signal input
rlabel metal2 s 46386 99200 46442 100000 6 wbd_adr_i[28]
port 42 nsew signal input
rlabel metal2 s 47398 99200 47454 100000 6 wbd_adr_i[29]
port 43 nsew signal input
rlabel metal2 s 20442 99200 20498 100000 6 wbd_adr_i[2]
port 44 nsew signal input
rlabel metal2 s 48410 99200 48466 100000 6 wbd_adr_i[30]
port 45 nsew signal input
rlabel metal2 s 49422 99200 49478 100000 6 wbd_adr_i[31]
port 46 nsew signal input
rlabel metal2 s 21454 99200 21510 100000 6 wbd_adr_i[3]
port 47 nsew signal input
rlabel metal2 s 22466 99200 22522 100000 6 wbd_adr_i[4]
port 48 nsew signal input
rlabel metal2 s 23386 99200 23442 100000 6 wbd_adr_i[5]
port 49 nsew signal input
rlabel metal2 s 24398 99200 24454 100000 6 wbd_adr_i[6]
port 50 nsew signal input
rlabel metal2 s 25410 99200 25466 100000 6 wbd_adr_i[7]
port 51 nsew signal input
rlabel metal2 s 26422 99200 26478 100000 6 wbd_adr_i[8]
port 52 nsew signal input
rlabel metal2 s 27434 99200 27490 100000 6 wbd_adr_i[9]
port 53 nsew signal input
rlabel metal2 s 54390 99200 54446 100000 6 wbd_dat_i[0]
port 54 nsew signal input
rlabel metal2 s 64418 99200 64474 100000 6 wbd_dat_i[10]
port 55 nsew signal input
rlabel metal2 s 65430 99200 65486 100000 6 wbd_dat_i[11]
port 56 nsew signal input
rlabel metal2 s 66442 99200 66498 100000 6 wbd_dat_i[12]
port 57 nsew signal input
rlabel metal2 s 67454 99200 67510 100000 6 wbd_dat_i[13]
port 58 nsew signal input
rlabel metal2 s 68374 99200 68430 100000 6 wbd_dat_i[14]
port 59 nsew signal input
rlabel metal2 s 69386 99200 69442 100000 6 wbd_dat_i[15]
port 60 nsew signal input
rlabel metal2 s 70398 99200 70454 100000 6 wbd_dat_i[16]
port 61 nsew signal input
rlabel metal2 s 71410 99200 71466 100000 6 wbd_dat_i[17]
port 62 nsew signal input
rlabel metal2 s 72422 99200 72478 100000 6 wbd_dat_i[18]
port 63 nsew signal input
rlabel metal2 s 73434 99200 73490 100000 6 wbd_dat_i[19]
port 64 nsew signal input
rlabel metal2 s 55402 99200 55458 100000 6 wbd_dat_i[1]
port 65 nsew signal input
rlabel metal2 s 74446 99200 74502 100000 6 wbd_dat_i[20]
port 66 nsew signal input
rlabel metal2 s 75458 99200 75514 100000 6 wbd_dat_i[21]
port 67 nsew signal input
rlabel metal2 s 76378 99200 76434 100000 6 wbd_dat_i[22]
port 68 nsew signal input
rlabel metal2 s 77390 99200 77446 100000 6 wbd_dat_i[23]
port 69 nsew signal input
rlabel metal2 s 78402 99200 78458 100000 6 wbd_dat_i[24]
port 70 nsew signal input
rlabel metal2 s 79414 99200 79470 100000 6 wbd_dat_i[25]
port 71 nsew signal input
rlabel metal2 s 80426 99200 80482 100000 6 wbd_dat_i[26]
port 72 nsew signal input
rlabel metal2 s 81438 99200 81494 100000 6 wbd_dat_i[27]
port 73 nsew signal input
rlabel metal2 s 82450 99200 82506 100000 6 wbd_dat_i[28]
port 74 nsew signal input
rlabel metal2 s 83370 99200 83426 100000 6 wbd_dat_i[29]
port 75 nsew signal input
rlabel metal2 s 56414 99200 56470 100000 6 wbd_dat_i[2]
port 76 nsew signal input
rlabel metal2 s 84382 99200 84438 100000 6 wbd_dat_i[30]
port 77 nsew signal input
rlabel metal2 s 85394 99200 85450 100000 6 wbd_dat_i[31]
port 78 nsew signal input
rlabel metal2 s 57426 99200 57482 100000 6 wbd_dat_i[3]
port 79 nsew signal input
rlabel metal2 s 58438 99200 58494 100000 6 wbd_dat_i[4]
port 80 nsew signal input
rlabel metal2 s 59450 99200 59506 100000 6 wbd_dat_i[5]
port 81 nsew signal input
rlabel metal2 s 60462 99200 60518 100000 6 wbd_dat_i[6]
port 82 nsew signal input
rlabel metal2 s 61382 99200 61438 100000 6 wbd_dat_i[7]
port 83 nsew signal input
rlabel metal2 s 62394 99200 62450 100000 6 wbd_dat_i[8]
port 84 nsew signal input
rlabel metal2 s 63406 99200 63462 100000 6 wbd_dat_i[9]
port 85 nsew signal input
rlabel metal2 s 86406 99200 86462 100000 6 wbd_dat_o[0]
port 86 nsew signal output
rlabel metal2 s 96434 99200 96490 100000 6 wbd_dat_o[10]
port 87 nsew signal output
rlabel metal2 s 97446 99200 97502 100000 6 wbd_dat_o[11]
port 88 nsew signal output
rlabel metal2 s 98366 99200 98422 100000 6 wbd_dat_o[12]
port 89 nsew signal output
rlabel metal2 s 99378 99200 99434 100000 6 wbd_dat_o[13]
port 90 nsew signal output
rlabel metal2 s 100390 99200 100446 100000 6 wbd_dat_o[14]
port 91 nsew signal output
rlabel metal2 s 101402 99200 101458 100000 6 wbd_dat_o[15]
port 92 nsew signal output
rlabel metal2 s 102414 99200 102470 100000 6 wbd_dat_o[16]
port 93 nsew signal output
rlabel metal2 s 103426 99200 103482 100000 6 wbd_dat_o[17]
port 94 nsew signal output
rlabel metal2 s 104438 99200 104494 100000 6 wbd_dat_o[18]
port 95 nsew signal output
rlabel metal2 s 105450 99200 105506 100000 6 wbd_dat_o[19]
port 96 nsew signal output
rlabel metal2 s 87418 99200 87474 100000 6 wbd_dat_o[1]
port 97 nsew signal output
rlabel metal2 s 106370 99200 106426 100000 6 wbd_dat_o[20]
port 98 nsew signal output
rlabel metal2 s 107382 99200 107438 100000 6 wbd_dat_o[21]
port 99 nsew signal output
rlabel metal2 s 108394 99200 108450 100000 6 wbd_dat_o[22]
port 100 nsew signal output
rlabel metal2 s 109406 99200 109462 100000 6 wbd_dat_o[23]
port 101 nsew signal output
rlabel metal2 s 110418 99200 110474 100000 6 wbd_dat_o[24]
port 102 nsew signal output
rlabel metal2 s 111430 99200 111486 100000 6 wbd_dat_o[25]
port 103 nsew signal output
rlabel metal2 s 112442 99200 112498 100000 6 wbd_dat_o[26]
port 104 nsew signal output
rlabel metal2 s 113362 99200 113418 100000 6 wbd_dat_o[27]
port 105 nsew signal output
rlabel metal2 s 114374 99200 114430 100000 6 wbd_dat_o[28]
port 106 nsew signal output
rlabel metal2 s 115386 99200 115442 100000 6 wbd_dat_o[29]
port 107 nsew signal output
rlabel metal2 s 88430 99200 88486 100000 6 wbd_dat_o[2]
port 108 nsew signal output
rlabel metal2 s 116398 99200 116454 100000 6 wbd_dat_o[30]
port 109 nsew signal output
rlabel metal2 s 117410 99200 117466 100000 6 wbd_dat_o[31]
port 110 nsew signal output
rlabel metal2 s 89442 99200 89498 100000 6 wbd_dat_o[3]
port 111 nsew signal output
rlabel metal2 s 90454 99200 90510 100000 6 wbd_dat_o[4]
port 112 nsew signal output
rlabel metal2 s 91374 99200 91430 100000 6 wbd_dat_o[5]
port 113 nsew signal output
rlabel metal2 s 92386 99200 92442 100000 6 wbd_dat_o[6]
port 114 nsew signal output
rlabel metal2 s 93398 99200 93454 100000 6 wbd_dat_o[7]
port 115 nsew signal output
rlabel metal2 s 94410 99200 94466 100000 6 wbd_dat_o[8]
port 116 nsew signal output
rlabel metal2 s 95422 99200 95478 100000 6 wbd_dat_o[9]
port 117 nsew signal output
rlabel metal2 s 119434 99200 119490 100000 6 wbd_err_o
port 118 nsew signal output
rlabel metal2 s 50434 99200 50490 100000 6 wbd_sel_i[0]
port 119 nsew signal input
rlabel metal2 s 51446 99200 51502 100000 6 wbd_sel_i[1]
port 120 nsew signal input
rlabel metal2 s 52458 99200 52514 100000 6 wbd_sel_i[2]
port 121 nsew signal input
rlabel metal2 s 53378 99200 53434 100000 6 wbd_sel_i[3]
port 122 nsew signal input
rlabel metal2 s 16394 99200 16450 100000 6 wbd_stb_i
port 123 nsew signal input
rlabel metal2 s 17406 99200 17462 100000 6 wbd_we_i
port 124 nsew signal input
rlabel metal4 s 96644 1040 96964 98512 6 VPWR
port 125 nsew power bidirectional
rlabel metal4 s 65924 1040 66244 98512 6 VPWR
port 126 nsew power bidirectional
rlabel metal4 s 35204 1040 35524 98512 6 VPWR
port 127 nsew power bidirectional
rlabel metal4 s 4484 1040 4804 98512 6 VPWR
port 128 nsew power bidirectional
rlabel metal5 s 1380 96118 118588 96438 6 VPWR
port 129 nsew power bidirectional
rlabel metal5 s 1380 65482 118588 65802 6 VPWR
port 130 nsew power bidirectional
rlabel metal5 s 1380 34846 118588 35166 6 VPWR
port 131 nsew power bidirectional
rlabel metal5 s 1380 4210 118588 4530 6 VPWR
port 132 nsew power bidirectional
rlabel metal4 s 112004 1040 112324 98512 6 VGND
port 133 nsew ground bidirectional
rlabel metal4 s 81284 1040 81604 98512 6 VGND
port 134 nsew ground bidirectional
rlabel metal4 s 50564 1040 50884 98512 6 VGND
port 135 nsew ground bidirectional
rlabel metal4 s 19844 1040 20164 98512 6 VGND
port 136 nsew ground bidirectional
rlabel metal5 s 1380 80800 118588 81120 6 VGND
port 137 nsew ground bidirectional
rlabel metal5 s 1380 50164 118588 50484 6 VGND
port 138 nsew ground bidirectional
rlabel metal5 s 1380 19528 118588 19848 6 VGND
port 139 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 120000 100000
string LEFview TRUE
string GDS_FILE /project/openlane/spi_master/runs/spi_master/results/magic/spim_top.gds
string GDS_END 10519404
string GDS_START 295934
<< end >>

