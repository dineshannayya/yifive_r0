magic
tech sky130A
magscale 1 2
timestamp 1623839057
<< obsli1 >>
rect 1104 2159 298816 237745
<< obsm1 >>
rect 750 1300 298816 237776
<< metal2 >>
rect 49974 239200 50030 240000
rect 149978 239200 150034 240000
rect 249982 239200 250038 240000
rect 754 0 810 800
rect 2226 0 2282 800
rect 3698 0 3754 800
rect 5170 0 5226 800
rect 6642 0 6698 800
rect 8114 0 8170 800
rect 9586 0 9642 800
rect 11058 0 11114 800
rect 12530 0 12586 800
rect 14002 0 14058 800
rect 15474 0 15530 800
rect 16946 0 17002 800
rect 18418 0 18474 800
rect 19890 0 19946 800
rect 21362 0 21418 800
rect 22834 0 22890 800
rect 24398 0 24454 800
rect 25870 0 25926 800
rect 27342 0 27398 800
rect 28814 0 28870 800
rect 30286 0 30342 800
rect 31758 0 31814 800
rect 33230 0 33286 800
rect 34702 0 34758 800
rect 36174 0 36230 800
rect 37646 0 37702 800
rect 39118 0 39174 800
rect 40590 0 40646 800
rect 42062 0 42118 800
rect 43534 0 43590 800
rect 45006 0 45062 800
rect 46478 0 46534 800
rect 48042 0 48098 800
rect 49514 0 49570 800
rect 50986 0 51042 800
rect 52458 0 52514 800
rect 53930 0 53986 800
rect 55402 0 55458 800
rect 56874 0 56930 800
rect 58346 0 58402 800
rect 59818 0 59874 800
rect 61290 0 61346 800
rect 62762 0 62818 800
rect 64234 0 64290 800
rect 65706 0 65762 800
rect 67178 0 67234 800
rect 68650 0 68706 800
rect 70214 0 70270 800
rect 71686 0 71742 800
rect 73158 0 73214 800
rect 74630 0 74686 800
rect 76102 0 76158 800
rect 77574 0 77630 800
rect 79046 0 79102 800
rect 80518 0 80574 800
rect 81990 0 82046 800
rect 83462 0 83518 800
rect 84934 0 84990 800
rect 86406 0 86462 800
rect 87878 0 87934 800
rect 89350 0 89406 800
rect 90822 0 90878 800
rect 92294 0 92350 800
rect 93858 0 93914 800
rect 95330 0 95386 800
rect 96802 0 96858 800
rect 98274 0 98330 800
rect 99746 0 99802 800
rect 101218 0 101274 800
rect 102690 0 102746 800
rect 104162 0 104218 800
rect 105634 0 105690 800
rect 107106 0 107162 800
rect 108578 0 108634 800
rect 110050 0 110106 800
rect 111522 0 111578 800
rect 112994 0 113050 800
rect 114466 0 114522 800
rect 115938 0 115994 800
rect 117502 0 117558 800
rect 118974 0 119030 800
rect 120446 0 120502 800
rect 121918 0 121974 800
rect 123390 0 123446 800
rect 124862 0 124918 800
rect 126334 0 126390 800
rect 127806 0 127862 800
rect 129278 0 129334 800
rect 130750 0 130806 800
rect 132222 0 132278 800
rect 133694 0 133750 800
rect 135166 0 135222 800
rect 136638 0 136694 800
rect 138110 0 138166 800
rect 139674 0 139730 800
rect 141146 0 141202 800
rect 142618 0 142674 800
rect 144090 0 144146 800
rect 145562 0 145618 800
rect 147034 0 147090 800
rect 148506 0 148562 800
rect 149978 0 150034 800
rect 151450 0 151506 800
rect 152922 0 152978 800
rect 154394 0 154450 800
rect 155866 0 155922 800
rect 157338 0 157394 800
rect 158810 0 158866 800
rect 160282 0 160338 800
rect 161754 0 161810 800
rect 163318 0 163374 800
rect 164790 0 164846 800
rect 166262 0 166318 800
rect 167734 0 167790 800
rect 169206 0 169262 800
rect 170678 0 170734 800
rect 172150 0 172206 800
rect 173622 0 173678 800
rect 175094 0 175150 800
rect 176566 0 176622 800
rect 178038 0 178094 800
rect 179510 0 179566 800
rect 180982 0 181038 800
rect 182454 0 182510 800
rect 183926 0 183982 800
rect 185490 0 185546 800
rect 186962 0 187018 800
rect 188434 0 188490 800
rect 189906 0 189962 800
rect 191378 0 191434 800
rect 192850 0 192906 800
rect 194322 0 194378 800
rect 195794 0 195850 800
rect 197266 0 197322 800
rect 198738 0 198794 800
rect 200210 0 200266 800
rect 201682 0 201738 800
rect 203154 0 203210 800
rect 204626 0 204682 800
rect 206098 0 206154 800
rect 207570 0 207626 800
rect 209134 0 209190 800
rect 210606 0 210662 800
rect 212078 0 212134 800
rect 213550 0 213606 800
rect 215022 0 215078 800
rect 216494 0 216550 800
rect 217966 0 218022 800
rect 219438 0 219494 800
rect 220910 0 220966 800
rect 222382 0 222438 800
rect 223854 0 223910 800
rect 225326 0 225382 800
rect 226798 0 226854 800
rect 228270 0 228326 800
rect 229742 0 229798 800
rect 231214 0 231270 800
rect 232778 0 232834 800
rect 234250 0 234306 800
rect 235722 0 235778 800
rect 237194 0 237250 800
rect 238666 0 238722 800
rect 240138 0 240194 800
rect 241610 0 241666 800
rect 243082 0 243138 800
rect 244554 0 244610 800
rect 246026 0 246082 800
rect 247498 0 247554 800
rect 248970 0 249026 800
rect 250442 0 250498 800
rect 251914 0 251970 800
rect 253386 0 253442 800
rect 254950 0 255006 800
rect 256422 0 256478 800
rect 257894 0 257950 800
rect 259366 0 259422 800
rect 260838 0 260894 800
rect 262310 0 262366 800
rect 263782 0 263838 800
rect 265254 0 265310 800
rect 266726 0 266782 800
rect 268198 0 268254 800
rect 269670 0 269726 800
rect 271142 0 271198 800
rect 272614 0 272670 800
rect 274086 0 274142 800
rect 275558 0 275614 800
rect 277030 0 277086 800
rect 278594 0 278650 800
rect 280066 0 280122 800
rect 281538 0 281594 800
rect 283010 0 283066 800
rect 284482 0 284538 800
rect 285954 0 286010 800
rect 287426 0 287482 800
rect 288898 0 288954 800
rect 290370 0 290426 800
rect 291842 0 291898 800
rect 293314 0 293370 800
rect 294786 0 294842 800
rect 296258 0 296314 800
rect 297730 0 297786 800
rect 299202 0 299258 800
<< obsm2 >>
rect 756 239144 49918 239200
rect 50086 239144 149922 239200
rect 150090 239144 249926 239200
rect 250094 239144 299258 239200
rect 756 856 299258 239144
rect 866 800 2170 856
rect 2338 800 3642 856
rect 3810 800 5114 856
rect 5282 800 6586 856
rect 6754 800 8058 856
rect 8226 800 9530 856
rect 9698 800 11002 856
rect 11170 800 12474 856
rect 12642 800 13946 856
rect 14114 800 15418 856
rect 15586 800 16890 856
rect 17058 800 18362 856
rect 18530 800 19834 856
rect 20002 800 21306 856
rect 21474 800 22778 856
rect 22946 800 24342 856
rect 24510 800 25814 856
rect 25982 800 27286 856
rect 27454 800 28758 856
rect 28926 800 30230 856
rect 30398 800 31702 856
rect 31870 800 33174 856
rect 33342 800 34646 856
rect 34814 800 36118 856
rect 36286 800 37590 856
rect 37758 800 39062 856
rect 39230 800 40534 856
rect 40702 800 42006 856
rect 42174 800 43478 856
rect 43646 800 44950 856
rect 45118 800 46422 856
rect 46590 800 47986 856
rect 48154 800 49458 856
rect 49626 800 50930 856
rect 51098 800 52402 856
rect 52570 800 53874 856
rect 54042 800 55346 856
rect 55514 800 56818 856
rect 56986 800 58290 856
rect 58458 800 59762 856
rect 59930 800 61234 856
rect 61402 800 62706 856
rect 62874 800 64178 856
rect 64346 800 65650 856
rect 65818 800 67122 856
rect 67290 800 68594 856
rect 68762 800 70158 856
rect 70326 800 71630 856
rect 71798 800 73102 856
rect 73270 800 74574 856
rect 74742 800 76046 856
rect 76214 800 77518 856
rect 77686 800 78990 856
rect 79158 800 80462 856
rect 80630 800 81934 856
rect 82102 800 83406 856
rect 83574 800 84878 856
rect 85046 800 86350 856
rect 86518 800 87822 856
rect 87990 800 89294 856
rect 89462 800 90766 856
rect 90934 800 92238 856
rect 92406 800 93802 856
rect 93970 800 95274 856
rect 95442 800 96746 856
rect 96914 800 98218 856
rect 98386 800 99690 856
rect 99858 800 101162 856
rect 101330 800 102634 856
rect 102802 800 104106 856
rect 104274 800 105578 856
rect 105746 800 107050 856
rect 107218 800 108522 856
rect 108690 800 109994 856
rect 110162 800 111466 856
rect 111634 800 112938 856
rect 113106 800 114410 856
rect 114578 800 115882 856
rect 116050 800 117446 856
rect 117614 800 118918 856
rect 119086 800 120390 856
rect 120558 800 121862 856
rect 122030 800 123334 856
rect 123502 800 124806 856
rect 124974 800 126278 856
rect 126446 800 127750 856
rect 127918 800 129222 856
rect 129390 800 130694 856
rect 130862 800 132166 856
rect 132334 800 133638 856
rect 133806 800 135110 856
rect 135278 800 136582 856
rect 136750 800 138054 856
rect 138222 800 139618 856
rect 139786 800 141090 856
rect 141258 800 142562 856
rect 142730 800 144034 856
rect 144202 800 145506 856
rect 145674 800 146978 856
rect 147146 800 148450 856
rect 148618 800 149922 856
rect 150090 800 151394 856
rect 151562 800 152866 856
rect 153034 800 154338 856
rect 154506 800 155810 856
rect 155978 800 157282 856
rect 157450 800 158754 856
rect 158922 800 160226 856
rect 160394 800 161698 856
rect 161866 800 163262 856
rect 163430 800 164734 856
rect 164902 800 166206 856
rect 166374 800 167678 856
rect 167846 800 169150 856
rect 169318 800 170622 856
rect 170790 800 172094 856
rect 172262 800 173566 856
rect 173734 800 175038 856
rect 175206 800 176510 856
rect 176678 800 177982 856
rect 178150 800 179454 856
rect 179622 800 180926 856
rect 181094 800 182398 856
rect 182566 800 183870 856
rect 184038 800 185434 856
rect 185602 800 186906 856
rect 187074 800 188378 856
rect 188546 800 189850 856
rect 190018 800 191322 856
rect 191490 800 192794 856
rect 192962 800 194266 856
rect 194434 800 195738 856
rect 195906 800 197210 856
rect 197378 800 198682 856
rect 198850 800 200154 856
rect 200322 800 201626 856
rect 201794 800 203098 856
rect 203266 800 204570 856
rect 204738 800 206042 856
rect 206210 800 207514 856
rect 207682 800 209078 856
rect 209246 800 210550 856
rect 210718 800 212022 856
rect 212190 800 213494 856
rect 213662 800 214966 856
rect 215134 800 216438 856
rect 216606 800 217910 856
rect 218078 800 219382 856
rect 219550 800 220854 856
rect 221022 800 222326 856
rect 222494 800 223798 856
rect 223966 800 225270 856
rect 225438 800 226742 856
rect 226910 800 228214 856
rect 228382 800 229686 856
rect 229854 800 231158 856
rect 231326 800 232722 856
rect 232890 800 234194 856
rect 234362 800 235666 856
rect 235834 800 237138 856
rect 237306 800 238610 856
rect 238778 800 240082 856
rect 240250 800 241554 856
rect 241722 800 243026 856
rect 243194 800 244498 856
rect 244666 800 245970 856
rect 246138 800 247442 856
rect 247610 800 248914 856
rect 249082 800 250386 856
rect 250554 800 251858 856
rect 252026 800 253330 856
rect 253498 800 254894 856
rect 255062 800 256366 856
rect 256534 800 257838 856
rect 258006 800 259310 856
rect 259478 800 260782 856
rect 260950 800 262254 856
rect 262422 800 263726 856
rect 263894 800 265198 856
rect 265366 800 266670 856
rect 266838 800 268142 856
rect 268310 800 269614 856
rect 269782 800 271086 856
rect 271254 800 272558 856
rect 272726 800 274030 856
rect 274198 800 275502 856
rect 275670 800 276974 856
rect 277142 800 278538 856
rect 278706 800 280010 856
rect 280178 800 281482 856
rect 281650 800 282954 856
rect 283122 800 284426 856
rect 284594 800 285898 856
rect 286066 800 287370 856
rect 287538 800 288842 856
rect 289010 800 290314 856
rect 290482 800 291786 856
rect 291954 800 293258 856
rect 293426 800 294730 856
rect 294898 800 296202 856
rect 296370 800 297674 856
rect 297842 800 299146 856
<< metal3 >>
rect 299200 237736 300000 237856
rect 299200 233384 300000 233504
rect 299200 229168 300000 229288
rect 299200 224816 300000 224936
rect 299200 220600 300000 220720
rect 299200 216248 300000 216368
rect 299200 212032 300000 212152
rect 299200 207680 300000 207800
rect 299200 203464 300000 203584
rect 299200 199112 300000 199232
rect 299200 194896 300000 195016
rect 299200 190544 300000 190664
rect 299200 186328 300000 186448
rect 299200 181976 300000 182096
rect 0 179936 800 180056
rect 299200 177760 300000 177880
rect 299200 173408 300000 173528
rect 299200 169192 300000 169312
rect 299200 164840 300000 164960
rect 299200 160624 300000 160744
rect 299200 156272 300000 156392
rect 299200 152056 300000 152176
rect 299200 147704 300000 147824
rect 299200 143488 300000 143608
rect 299200 139136 300000 139256
rect 299200 134920 300000 135040
rect 299200 130568 300000 130688
rect 299200 126352 300000 126472
rect 299200 122000 300000 122120
rect 299200 117648 300000 117768
rect 299200 113432 300000 113552
rect 299200 109080 300000 109200
rect 299200 104864 300000 104984
rect 299200 100512 300000 100632
rect 299200 96296 300000 96416
rect 299200 91944 300000 92064
rect 299200 87728 300000 87848
rect 299200 83376 300000 83496
rect 299200 79160 300000 79280
rect 299200 74808 300000 74928
rect 299200 70592 300000 70712
rect 299200 66240 300000 66360
rect 299200 62024 300000 62144
rect 0 59984 800 60104
rect 299200 57672 300000 57792
rect 299200 53456 300000 53576
rect 299200 49104 300000 49224
rect 299200 44888 300000 45008
rect 299200 40536 300000 40656
rect 299200 36320 300000 36440
rect 299200 31968 300000 32088
rect 299200 27752 300000 27872
rect 299200 23400 300000 23520
rect 299200 19184 300000 19304
rect 299200 14832 300000 14952
rect 299200 10616 300000 10736
rect 299200 6264 300000 6384
rect 299200 2048 300000 2168
<< obsm3 >>
rect 800 237656 299120 237829
rect 800 233584 299263 237656
rect 800 233304 299120 233584
rect 800 229368 299263 233304
rect 800 229088 299120 229368
rect 800 225016 299263 229088
rect 800 224736 299120 225016
rect 800 220800 299263 224736
rect 800 220520 299120 220800
rect 800 216448 299263 220520
rect 800 216168 299120 216448
rect 800 212232 299263 216168
rect 800 211952 299120 212232
rect 800 207880 299263 211952
rect 800 207600 299120 207880
rect 800 203664 299263 207600
rect 800 203384 299120 203664
rect 800 199312 299263 203384
rect 800 199032 299120 199312
rect 800 195096 299263 199032
rect 800 194816 299120 195096
rect 800 190744 299263 194816
rect 800 190464 299120 190744
rect 800 186528 299263 190464
rect 800 186248 299120 186528
rect 800 182176 299263 186248
rect 800 181896 299120 182176
rect 800 180136 299263 181896
rect 880 179856 299263 180136
rect 800 177960 299263 179856
rect 800 177680 299120 177960
rect 800 173608 299263 177680
rect 800 173328 299120 173608
rect 800 169392 299263 173328
rect 800 169112 299120 169392
rect 800 165040 299263 169112
rect 800 164760 299120 165040
rect 800 160824 299263 164760
rect 800 160544 299120 160824
rect 800 156472 299263 160544
rect 800 156192 299120 156472
rect 800 152256 299263 156192
rect 800 151976 299120 152256
rect 800 147904 299263 151976
rect 800 147624 299120 147904
rect 800 143688 299263 147624
rect 800 143408 299120 143688
rect 800 139336 299263 143408
rect 800 139056 299120 139336
rect 800 135120 299263 139056
rect 800 134840 299120 135120
rect 800 130768 299263 134840
rect 800 130488 299120 130768
rect 800 126552 299263 130488
rect 800 126272 299120 126552
rect 800 122200 299263 126272
rect 800 121920 299120 122200
rect 800 117848 299263 121920
rect 800 117568 299120 117848
rect 800 113632 299263 117568
rect 800 113352 299120 113632
rect 800 109280 299263 113352
rect 800 109000 299120 109280
rect 800 105064 299263 109000
rect 800 104784 299120 105064
rect 800 100712 299263 104784
rect 800 100432 299120 100712
rect 800 96496 299263 100432
rect 800 96216 299120 96496
rect 800 92144 299263 96216
rect 800 91864 299120 92144
rect 800 87928 299263 91864
rect 800 87648 299120 87928
rect 800 83576 299263 87648
rect 800 83296 299120 83576
rect 800 79360 299263 83296
rect 800 79080 299120 79360
rect 800 75008 299263 79080
rect 800 74728 299120 75008
rect 800 70792 299263 74728
rect 800 70512 299120 70792
rect 800 66440 299263 70512
rect 800 66160 299120 66440
rect 800 62224 299263 66160
rect 800 61944 299120 62224
rect 800 60184 299263 61944
rect 880 59904 299263 60184
rect 800 57872 299263 59904
rect 800 57592 299120 57872
rect 800 53656 299263 57592
rect 800 53376 299120 53656
rect 800 49304 299263 53376
rect 800 49024 299120 49304
rect 800 45088 299263 49024
rect 800 44808 299120 45088
rect 800 40736 299263 44808
rect 800 40456 299120 40736
rect 800 36520 299263 40456
rect 800 36240 299120 36520
rect 800 32168 299263 36240
rect 800 31888 299120 32168
rect 800 27952 299263 31888
rect 800 27672 299120 27952
rect 800 23600 299263 27672
rect 800 23320 299120 23600
rect 800 19384 299263 23320
rect 800 19104 299120 19384
rect 800 15032 299263 19104
rect 800 14752 299120 15032
rect 800 10816 299263 14752
rect 800 10536 299120 10816
rect 800 6464 299263 10536
rect 800 6184 299120 6464
rect 800 2248 299263 6184
rect 800 2075 299120 2248
<< metal4 >>
rect 4208 2128 4528 237776
rect 19568 2128 19888 237776
rect 34928 2128 35248 237776
rect 50288 2128 50608 237776
rect 65648 2128 65968 237776
rect 81008 2128 81328 237776
rect 96368 2128 96688 237776
rect 111728 2128 112048 237776
rect 127088 2128 127408 237776
rect 142448 2128 142768 237776
rect 157808 2128 158128 237776
rect 173168 2128 173488 237776
rect 188528 2128 188848 237776
rect 203888 2128 204208 237776
rect 219248 2128 219568 237776
rect 234608 2128 234928 237776
rect 249968 2128 250288 237776
rect 265328 2128 265648 237776
rect 280688 2128 281008 237776
rect 296048 2128 296368 237776
<< obsm4 >>
rect 65379 11731 65568 156365
rect 66048 11731 80928 156365
rect 81408 11731 96288 156365
rect 96768 11731 111648 156365
rect 112128 11731 127008 156365
rect 127488 11731 142368 156365
rect 142848 11731 157728 156365
rect 158208 11731 173088 156365
rect 173568 11731 188448 156365
rect 188928 11731 203808 156365
rect 204288 11731 219168 156365
rect 219648 11731 234528 156365
rect 235008 11731 241717 156365
<< metal5 >>
rect 1104 235068 298816 235388
rect 1104 219750 298816 220070
rect 1104 204432 298816 204752
rect 1104 189114 298816 189434
rect 1104 173796 298816 174116
rect 1104 158478 298816 158798
rect 1104 143160 298816 143480
rect 1104 127842 298816 128162
rect 1104 112524 298816 112844
rect 1104 97206 298816 97526
rect 1104 81888 298816 82208
rect 1104 66570 298816 66890
rect 1104 51252 298816 51572
rect 1104 35934 298816 36254
rect 1104 20616 298816 20936
rect 1104 5298 298816 5618
<< labels >>
rlabel metal3 s 299200 2048 300000 2168 6 clk
port 1 nsew signal input
rlabel metal3 s 299200 6264 300000 6384 6 cpu_rst_n
port 2 nsew signal input
rlabel metal3 s 299200 96296 300000 96416 6 fuse_mhartid[0]
port 3 nsew signal input
rlabel metal3 s 299200 139136 300000 139256 6 fuse_mhartid[10]
port 4 nsew signal input
rlabel metal3 s 299200 143488 300000 143608 6 fuse_mhartid[11]
port 5 nsew signal input
rlabel metal3 s 299200 147704 300000 147824 6 fuse_mhartid[12]
port 6 nsew signal input
rlabel metal3 s 299200 152056 300000 152176 6 fuse_mhartid[13]
port 7 nsew signal input
rlabel metal3 s 299200 156272 300000 156392 6 fuse_mhartid[14]
port 8 nsew signal input
rlabel metal3 s 299200 160624 300000 160744 6 fuse_mhartid[15]
port 9 nsew signal input
rlabel metal3 s 299200 164840 300000 164960 6 fuse_mhartid[16]
port 10 nsew signal input
rlabel metal3 s 299200 169192 300000 169312 6 fuse_mhartid[17]
port 11 nsew signal input
rlabel metal3 s 299200 173408 300000 173528 6 fuse_mhartid[18]
port 12 nsew signal input
rlabel metal3 s 299200 177760 300000 177880 6 fuse_mhartid[19]
port 13 nsew signal input
rlabel metal3 s 299200 100512 300000 100632 6 fuse_mhartid[1]
port 14 nsew signal input
rlabel metal3 s 299200 181976 300000 182096 6 fuse_mhartid[20]
port 15 nsew signal input
rlabel metal3 s 299200 186328 300000 186448 6 fuse_mhartid[21]
port 16 nsew signal input
rlabel metal3 s 299200 190544 300000 190664 6 fuse_mhartid[22]
port 17 nsew signal input
rlabel metal3 s 299200 194896 300000 195016 6 fuse_mhartid[23]
port 18 nsew signal input
rlabel metal3 s 299200 199112 300000 199232 6 fuse_mhartid[24]
port 19 nsew signal input
rlabel metal3 s 299200 203464 300000 203584 6 fuse_mhartid[25]
port 20 nsew signal input
rlabel metal3 s 299200 207680 300000 207800 6 fuse_mhartid[26]
port 21 nsew signal input
rlabel metal3 s 299200 212032 300000 212152 6 fuse_mhartid[27]
port 22 nsew signal input
rlabel metal3 s 299200 216248 300000 216368 6 fuse_mhartid[28]
port 23 nsew signal input
rlabel metal3 s 299200 220600 300000 220720 6 fuse_mhartid[29]
port 24 nsew signal input
rlabel metal3 s 299200 104864 300000 104984 6 fuse_mhartid[2]
port 25 nsew signal input
rlabel metal3 s 299200 224816 300000 224936 6 fuse_mhartid[30]
port 26 nsew signal input
rlabel metal3 s 299200 229168 300000 229288 6 fuse_mhartid[31]
port 27 nsew signal input
rlabel metal3 s 299200 109080 300000 109200 6 fuse_mhartid[3]
port 28 nsew signal input
rlabel metal3 s 299200 113432 300000 113552 6 fuse_mhartid[4]
port 29 nsew signal input
rlabel metal3 s 299200 117648 300000 117768 6 fuse_mhartid[5]
port 30 nsew signal input
rlabel metal3 s 299200 122000 300000 122120 6 fuse_mhartid[6]
port 31 nsew signal input
rlabel metal3 s 299200 126352 300000 126472 6 fuse_mhartid[7]
port 32 nsew signal input
rlabel metal3 s 299200 130568 300000 130688 6 fuse_mhartid[8]
port 33 nsew signal input
rlabel metal3 s 299200 134920 300000 135040 6 fuse_mhartid[9]
port 34 nsew signal input
rlabel metal3 s 299200 10616 300000 10736 6 irq_lines[0]
port 35 nsew signal input
rlabel metal3 s 299200 53456 300000 53576 6 irq_lines[10]
port 36 nsew signal input
rlabel metal3 s 299200 57672 300000 57792 6 irq_lines[11]
port 37 nsew signal input
rlabel metal3 s 299200 62024 300000 62144 6 irq_lines[12]
port 38 nsew signal input
rlabel metal3 s 299200 66240 300000 66360 6 irq_lines[13]
port 39 nsew signal input
rlabel metal3 s 299200 70592 300000 70712 6 irq_lines[14]
port 40 nsew signal input
rlabel metal3 s 299200 74808 300000 74928 6 irq_lines[15]
port 41 nsew signal input
rlabel metal3 s 299200 14832 300000 14952 6 irq_lines[1]
port 42 nsew signal input
rlabel metal3 s 299200 19184 300000 19304 6 irq_lines[2]
port 43 nsew signal input
rlabel metal3 s 299200 23400 300000 23520 6 irq_lines[3]
port 44 nsew signal input
rlabel metal3 s 299200 27752 300000 27872 6 irq_lines[4]
port 45 nsew signal input
rlabel metal3 s 299200 31968 300000 32088 6 irq_lines[5]
port 46 nsew signal input
rlabel metal3 s 299200 36320 300000 36440 6 irq_lines[6]
port 47 nsew signal input
rlabel metal3 s 299200 40536 300000 40656 6 irq_lines[7]
port 48 nsew signal input
rlabel metal3 s 299200 44888 300000 45008 6 irq_lines[8]
port 49 nsew signal input
rlabel metal3 s 299200 49104 300000 49224 6 irq_lines[9]
port 50 nsew signal input
rlabel metal3 s 299200 79160 300000 79280 6 pwrup_rst_n
port 51 nsew signal input
rlabel metal3 s 299200 83376 300000 83496 6 rst_n
port 52 nsew signal input
rlabel metal3 s 299200 87728 300000 87848 6 rtc_clk
port 53 nsew signal input
rlabel metal3 s 299200 91944 300000 92064 6 soft_irq
port 54 nsew signal input
rlabel metal3 s 0 59984 800 60104 6 test_mode
port 55 nsew signal input
rlabel metal3 s 0 179936 800 180056 6 test_rst_n
port 56 nsew signal input
rlabel metal2 s 293314 0 293370 800 6 wbd_dmem_ack_i
port 57 nsew signal input
rlabel metal2 s 149978 0 150034 800 6 wbd_dmem_adr_o[0]
port 58 nsew signal output
rlabel metal2 s 164790 0 164846 800 6 wbd_dmem_adr_o[10]
port 59 nsew signal output
rlabel metal2 s 166262 0 166318 800 6 wbd_dmem_adr_o[11]
port 60 nsew signal output
rlabel metal2 s 167734 0 167790 800 6 wbd_dmem_adr_o[12]
port 61 nsew signal output
rlabel metal2 s 169206 0 169262 800 6 wbd_dmem_adr_o[13]
port 62 nsew signal output
rlabel metal2 s 170678 0 170734 800 6 wbd_dmem_adr_o[14]
port 63 nsew signal output
rlabel metal2 s 172150 0 172206 800 6 wbd_dmem_adr_o[15]
port 64 nsew signal output
rlabel metal2 s 173622 0 173678 800 6 wbd_dmem_adr_o[16]
port 65 nsew signal output
rlabel metal2 s 175094 0 175150 800 6 wbd_dmem_adr_o[17]
port 66 nsew signal output
rlabel metal2 s 176566 0 176622 800 6 wbd_dmem_adr_o[18]
port 67 nsew signal output
rlabel metal2 s 178038 0 178094 800 6 wbd_dmem_adr_o[19]
port 68 nsew signal output
rlabel metal2 s 151450 0 151506 800 6 wbd_dmem_adr_o[1]
port 69 nsew signal output
rlabel metal2 s 179510 0 179566 800 6 wbd_dmem_adr_o[20]
port 70 nsew signal output
rlabel metal2 s 180982 0 181038 800 6 wbd_dmem_adr_o[21]
port 71 nsew signal output
rlabel metal2 s 182454 0 182510 800 6 wbd_dmem_adr_o[22]
port 72 nsew signal output
rlabel metal2 s 183926 0 183982 800 6 wbd_dmem_adr_o[23]
port 73 nsew signal output
rlabel metal2 s 185490 0 185546 800 6 wbd_dmem_adr_o[24]
port 74 nsew signal output
rlabel metal2 s 186962 0 187018 800 6 wbd_dmem_adr_o[25]
port 75 nsew signal output
rlabel metal2 s 188434 0 188490 800 6 wbd_dmem_adr_o[26]
port 76 nsew signal output
rlabel metal2 s 189906 0 189962 800 6 wbd_dmem_adr_o[27]
port 77 nsew signal output
rlabel metal2 s 191378 0 191434 800 6 wbd_dmem_adr_o[28]
port 78 nsew signal output
rlabel metal2 s 192850 0 192906 800 6 wbd_dmem_adr_o[29]
port 79 nsew signal output
rlabel metal2 s 152922 0 152978 800 6 wbd_dmem_adr_o[2]
port 80 nsew signal output
rlabel metal2 s 194322 0 194378 800 6 wbd_dmem_adr_o[30]
port 81 nsew signal output
rlabel metal2 s 195794 0 195850 800 6 wbd_dmem_adr_o[31]
port 82 nsew signal output
rlabel metal2 s 154394 0 154450 800 6 wbd_dmem_adr_o[3]
port 83 nsew signal output
rlabel metal2 s 155866 0 155922 800 6 wbd_dmem_adr_o[4]
port 84 nsew signal output
rlabel metal2 s 157338 0 157394 800 6 wbd_dmem_adr_o[5]
port 85 nsew signal output
rlabel metal2 s 158810 0 158866 800 6 wbd_dmem_adr_o[6]
port 86 nsew signal output
rlabel metal2 s 160282 0 160338 800 6 wbd_dmem_adr_o[7]
port 87 nsew signal output
rlabel metal2 s 161754 0 161810 800 6 wbd_dmem_adr_o[8]
port 88 nsew signal output
rlabel metal2 s 163318 0 163374 800 6 wbd_dmem_adr_o[9]
port 89 nsew signal output
rlabel metal2 s 246026 0 246082 800 6 wbd_dmem_dat_i[0]
port 90 nsew signal input
rlabel metal2 s 260838 0 260894 800 6 wbd_dmem_dat_i[10]
port 91 nsew signal input
rlabel metal2 s 262310 0 262366 800 6 wbd_dmem_dat_i[11]
port 92 nsew signal input
rlabel metal2 s 263782 0 263838 800 6 wbd_dmem_dat_i[12]
port 93 nsew signal input
rlabel metal2 s 265254 0 265310 800 6 wbd_dmem_dat_i[13]
port 94 nsew signal input
rlabel metal2 s 266726 0 266782 800 6 wbd_dmem_dat_i[14]
port 95 nsew signal input
rlabel metal2 s 268198 0 268254 800 6 wbd_dmem_dat_i[15]
port 96 nsew signal input
rlabel metal2 s 269670 0 269726 800 6 wbd_dmem_dat_i[16]
port 97 nsew signal input
rlabel metal2 s 271142 0 271198 800 6 wbd_dmem_dat_i[17]
port 98 nsew signal input
rlabel metal2 s 272614 0 272670 800 6 wbd_dmem_dat_i[18]
port 99 nsew signal input
rlabel metal2 s 274086 0 274142 800 6 wbd_dmem_dat_i[19]
port 100 nsew signal input
rlabel metal2 s 247498 0 247554 800 6 wbd_dmem_dat_i[1]
port 101 nsew signal input
rlabel metal2 s 275558 0 275614 800 6 wbd_dmem_dat_i[20]
port 102 nsew signal input
rlabel metal2 s 277030 0 277086 800 6 wbd_dmem_dat_i[21]
port 103 nsew signal input
rlabel metal2 s 278594 0 278650 800 6 wbd_dmem_dat_i[22]
port 104 nsew signal input
rlabel metal2 s 280066 0 280122 800 6 wbd_dmem_dat_i[23]
port 105 nsew signal input
rlabel metal2 s 281538 0 281594 800 6 wbd_dmem_dat_i[24]
port 106 nsew signal input
rlabel metal2 s 283010 0 283066 800 6 wbd_dmem_dat_i[25]
port 107 nsew signal input
rlabel metal2 s 284482 0 284538 800 6 wbd_dmem_dat_i[26]
port 108 nsew signal input
rlabel metal2 s 285954 0 286010 800 6 wbd_dmem_dat_i[27]
port 109 nsew signal input
rlabel metal2 s 287426 0 287482 800 6 wbd_dmem_dat_i[28]
port 110 nsew signal input
rlabel metal2 s 288898 0 288954 800 6 wbd_dmem_dat_i[29]
port 111 nsew signal input
rlabel metal2 s 248970 0 249026 800 6 wbd_dmem_dat_i[2]
port 112 nsew signal input
rlabel metal2 s 290370 0 290426 800 6 wbd_dmem_dat_i[30]
port 113 nsew signal input
rlabel metal2 s 291842 0 291898 800 6 wbd_dmem_dat_i[31]
port 114 nsew signal input
rlabel metal2 s 250442 0 250498 800 6 wbd_dmem_dat_i[3]
port 115 nsew signal input
rlabel metal2 s 251914 0 251970 800 6 wbd_dmem_dat_i[4]
port 116 nsew signal input
rlabel metal2 s 253386 0 253442 800 6 wbd_dmem_dat_i[5]
port 117 nsew signal input
rlabel metal2 s 254950 0 255006 800 6 wbd_dmem_dat_i[6]
port 118 nsew signal input
rlabel metal2 s 256422 0 256478 800 6 wbd_dmem_dat_i[7]
port 119 nsew signal input
rlabel metal2 s 257894 0 257950 800 6 wbd_dmem_dat_i[8]
port 120 nsew signal input
rlabel metal2 s 259366 0 259422 800 6 wbd_dmem_dat_i[9]
port 121 nsew signal input
rlabel metal2 s 198738 0 198794 800 6 wbd_dmem_dat_o[0]
port 122 nsew signal output
rlabel metal2 s 213550 0 213606 800 6 wbd_dmem_dat_o[10]
port 123 nsew signal output
rlabel metal2 s 215022 0 215078 800 6 wbd_dmem_dat_o[11]
port 124 nsew signal output
rlabel metal2 s 216494 0 216550 800 6 wbd_dmem_dat_o[12]
port 125 nsew signal output
rlabel metal2 s 217966 0 218022 800 6 wbd_dmem_dat_o[13]
port 126 nsew signal output
rlabel metal2 s 219438 0 219494 800 6 wbd_dmem_dat_o[14]
port 127 nsew signal output
rlabel metal2 s 220910 0 220966 800 6 wbd_dmem_dat_o[15]
port 128 nsew signal output
rlabel metal2 s 222382 0 222438 800 6 wbd_dmem_dat_o[16]
port 129 nsew signal output
rlabel metal2 s 223854 0 223910 800 6 wbd_dmem_dat_o[17]
port 130 nsew signal output
rlabel metal2 s 225326 0 225382 800 6 wbd_dmem_dat_o[18]
port 131 nsew signal output
rlabel metal2 s 226798 0 226854 800 6 wbd_dmem_dat_o[19]
port 132 nsew signal output
rlabel metal2 s 200210 0 200266 800 6 wbd_dmem_dat_o[1]
port 133 nsew signal output
rlabel metal2 s 228270 0 228326 800 6 wbd_dmem_dat_o[20]
port 134 nsew signal output
rlabel metal2 s 229742 0 229798 800 6 wbd_dmem_dat_o[21]
port 135 nsew signal output
rlabel metal2 s 231214 0 231270 800 6 wbd_dmem_dat_o[22]
port 136 nsew signal output
rlabel metal2 s 232778 0 232834 800 6 wbd_dmem_dat_o[23]
port 137 nsew signal output
rlabel metal2 s 234250 0 234306 800 6 wbd_dmem_dat_o[24]
port 138 nsew signal output
rlabel metal2 s 235722 0 235778 800 6 wbd_dmem_dat_o[25]
port 139 nsew signal output
rlabel metal2 s 237194 0 237250 800 6 wbd_dmem_dat_o[26]
port 140 nsew signal output
rlabel metal2 s 238666 0 238722 800 6 wbd_dmem_dat_o[27]
port 141 nsew signal output
rlabel metal2 s 240138 0 240194 800 6 wbd_dmem_dat_o[28]
port 142 nsew signal output
rlabel metal2 s 241610 0 241666 800 6 wbd_dmem_dat_o[29]
port 143 nsew signal output
rlabel metal2 s 201682 0 201738 800 6 wbd_dmem_dat_o[2]
port 144 nsew signal output
rlabel metal2 s 243082 0 243138 800 6 wbd_dmem_dat_o[30]
port 145 nsew signal output
rlabel metal2 s 244554 0 244610 800 6 wbd_dmem_dat_o[31]
port 146 nsew signal output
rlabel metal2 s 203154 0 203210 800 6 wbd_dmem_dat_o[3]
port 147 nsew signal output
rlabel metal2 s 204626 0 204682 800 6 wbd_dmem_dat_o[4]
port 148 nsew signal output
rlabel metal2 s 206098 0 206154 800 6 wbd_dmem_dat_o[5]
port 149 nsew signal output
rlabel metal2 s 207570 0 207626 800 6 wbd_dmem_dat_o[6]
port 150 nsew signal output
rlabel metal2 s 209134 0 209190 800 6 wbd_dmem_dat_o[7]
port 151 nsew signal output
rlabel metal2 s 210606 0 210662 800 6 wbd_dmem_dat_o[8]
port 152 nsew signal output
rlabel metal2 s 212078 0 212134 800 6 wbd_dmem_dat_o[9]
port 153 nsew signal output
rlabel metal2 s 294786 0 294842 800 6 wbd_dmem_err_i
port 154 nsew signal input
rlabel metal2 s 296258 0 296314 800 6 wbd_dmem_sel_o[0]
port 155 nsew signal output
rlabel metal2 s 49974 239200 50030 240000 6 wbd_dmem_sel_o[1]
port 156 nsew signal output
rlabel metal3 s 299200 237736 300000 237856 6 wbd_dmem_sel_o[2]
port 157 nsew signal output
rlabel metal2 s 299202 0 299258 800 6 wbd_dmem_sel_o[3]
port 158 nsew signal output
rlabel metal2 s 148506 0 148562 800 6 wbd_dmem_stb_o
port 159 nsew signal output
rlabel metal2 s 197266 0 197322 800 6 wbd_dmem_we_o
port 160 nsew signal output
rlabel metal2 s 145562 0 145618 800 6 wbd_imem_ack_i
port 161 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbd_imem_adr_o[0]
port 162 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 wbd_imem_adr_o[10]
port 163 nsew signal output
rlabel metal2 s 19890 0 19946 800 6 wbd_imem_adr_o[11]
port 164 nsew signal output
rlabel metal2 s 21362 0 21418 800 6 wbd_imem_adr_o[12]
port 165 nsew signal output
rlabel metal2 s 22834 0 22890 800 6 wbd_imem_adr_o[13]
port 166 nsew signal output
rlabel metal2 s 24398 0 24454 800 6 wbd_imem_adr_o[14]
port 167 nsew signal output
rlabel metal2 s 25870 0 25926 800 6 wbd_imem_adr_o[15]
port 168 nsew signal output
rlabel metal2 s 27342 0 27398 800 6 wbd_imem_adr_o[16]
port 169 nsew signal output
rlabel metal2 s 28814 0 28870 800 6 wbd_imem_adr_o[17]
port 170 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 wbd_imem_adr_o[18]
port 171 nsew signal output
rlabel metal2 s 31758 0 31814 800 6 wbd_imem_adr_o[19]
port 172 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 wbd_imem_adr_o[1]
port 173 nsew signal output
rlabel metal2 s 33230 0 33286 800 6 wbd_imem_adr_o[20]
port 174 nsew signal output
rlabel metal2 s 34702 0 34758 800 6 wbd_imem_adr_o[21]
port 175 nsew signal output
rlabel metal2 s 36174 0 36230 800 6 wbd_imem_adr_o[22]
port 176 nsew signal output
rlabel metal2 s 37646 0 37702 800 6 wbd_imem_adr_o[23]
port 177 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 wbd_imem_adr_o[24]
port 178 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 wbd_imem_adr_o[25]
port 179 nsew signal output
rlabel metal2 s 42062 0 42118 800 6 wbd_imem_adr_o[26]
port 180 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 wbd_imem_adr_o[27]
port 181 nsew signal output
rlabel metal2 s 45006 0 45062 800 6 wbd_imem_adr_o[28]
port 182 nsew signal output
rlabel metal2 s 46478 0 46534 800 6 wbd_imem_adr_o[29]
port 183 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 wbd_imem_adr_o[2]
port 184 nsew signal output
rlabel metal2 s 48042 0 48098 800 6 wbd_imem_adr_o[30]
port 185 nsew signal output
rlabel metal2 s 49514 0 49570 800 6 wbd_imem_adr_o[31]
port 186 nsew signal output
rlabel metal2 s 8114 0 8170 800 6 wbd_imem_adr_o[3]
port 187 nsew signal output
rlabel metal2 s 9586 0 9642 800 6 wbd_imem_adr_o[4]
port 188 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 wbd_imem_adr_o[5]
port 189 nsew signal output
rlabel metal2 s 12530 0 12586 800 6 wbd_imem_adr_o[6]
port 190 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 wbd_imem_adr_o[7]
port 191 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 wbd_imem_adr_o[8]
port 192 nsew signal output
rlabel metal2 s 16946 0 17002 800 6 wbd_imem_adr_o[9]
port 193 nsew signal output
rlabel metal2 s 98274 0 98330 800 6 wbd_imem_dat_i[0]
port 194 nsew signal input
rlabel metal2 s 112994 0 113050 800 6 wbd_imem_dat_i[10]
port 195 nsew signal input
rlabel metal2 s 114466 0 114522 800 6 wbd_imem_dat_i[11]
port 196 nsew signal input
rlabel metal2 s 115938 0 115994 800 6 wbd_imem_dat_i[12]
port 197 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 wbd_imem_dat_i[13]
port 198 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 wbd_imem_dat_i[14]
port 199 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 wbd_imem_dat_i[15]
port 200 nsew signal input
rlabel metal2 s 121918 0 121974 800 6 wbd_imem_dat_i[16]
port 201 nsew signal input
rlabel metal2 s 123390 0 123446 800 6 wbd_imem_dat_i[17]
port 202 nsew signal input
rlabel metal2 s 124862 0 124918 800 6 wbd_imem_dat_i[18]
port 203 nsew signal input
rlabel metal2 s 126334 0 126390 800 6 wbd_imem_dat_i[19]
port 204 nsew signal input
rlabel metal2 s 99746 0 99802 800 6 wbd_imem_dat_i[1]
port 205 nsew signal input
rlabel metal2 s 127806 0 127862 800 6 wbd_imem_dat_i[20]
port 206 nsew signal input
rlabel metal2 s 129278 0 129334 800 6 wbd_imem_dat_i[21]
port 207 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 wbd_imem_dat_i[22]
port 208 nsew signal input
rlabel metal2 s 132222 0 132278 800 6 wbd_imem_dat_i[23]
port 209 nsew signal input
rlabel metal2 s 133694 0 133750 800 6 wbd_imem_dat_i[24]
port 210 nsew signal input
rlabel metal2 s 135166 0 135222 800 6 wbd_imem_dat_i[25]
port 211 nsew signal input
rlabel metal2 s 136638 0 136694 800 6 wbd_imem_dat_i[26]
port 212 nsew signal input
rlabel metal2 s 138110 0 138166 800 6 wbd_imem_dat_i[27]
port 213 nsew signal input
rlabel metal2 s 139674 0 139730 800 6 wbd_imem_dat_i[28]
port 214 nsew signal input
rlabel metal2 s 141146 0 141202 800 6 wbd_imem_dat_i[29]
port 215 nsew signal input
rlabel metal2 s 101218 0 101274 800 6 wbd_imem_dat_i[2]
port 216 nsew signal input
rlabel metal2 s 142618 0 142674 800 6 wbd_imem_dat_i[30]
port 217 nsew signal input
rlabel metal2 s 144090 0 144146 800 6 wbd_imem_dat_i[31]
port 218 nsew signal input
rlabel metal2 s 102690 0 102746 800 6 wbd_imem_dat_i[3]
port 219 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 wbd_imem_dat_i[4]
port 220 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 wbd_imem_dat_i[5]
port 221 nsew signal input
rlabel metal2 s 107106 0 107162 800 6 wbd_imem_dat_i[6]
port 222 nsew signal input
rlabel metal2 s 108578 0 108634 800 6 wbd_imem_dat_i[7]
port 223 nsew signal input
rlabel metal2 s 110050 0 110106 800 6 wbd_imem_dat_i[8]
port 224 nsew signal input
rlabel metal2 s 111522 0 111578 800 6 wbd_imem_dat_i[9]
port 225 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 wbd_imem_dat_o[0]
port 226 nsew signal output
rlabel metal2 s 65706 0 65762 800 6 wbd_imem_dat_o[10]
port 227 nsew signal output
rlabel metal2 s 67178 0 67234 800 6 wbd_imem_dat_o[11]
port 228 nsew signal output
rlabel metal2 s 68650 0 68706 800 6 wbd_imem_dat_o[12]
port 229 nsew signal output
rlabel metal2 s 70214 0 70270 800 6 wbd_imem_dat_o[13]
port 230 nsew signal output
rlabel metal2 s 71686 0 71742 800 6 wbd_imem_dat_o[14]
port 231 nsew signal output
rlabel metal2 s 73158 0 73214 800 6 wbd_imem_dat_o[15]
port 232 nsew signal output
rlabel metal2 s 74630 0 74686 800 6 wbd_imem_dat_o[16]
port 233 nsew signal output
rlabel metal2 s 76102 0 76158 800 6 wbd_imem_dat_o[17]
port 234 nsew signal output
rlabel metal2 s 77574 0 77630 800 6 wbd_imem_dat_o[18]
port 235 nsew signal output
rlabel metal2 s 79046 0 79102 800 6 wbd_imem_dat_o[19]
port 236 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 wbd_imem_dat_o[1]
port 237 nsew signal output
rlabel metal2 s 80518 0 80574 800 6 wbd_imem_dat_o[20]
port 238 nsew signal output
rlabel metal2 s 81990 0 82046 800 6 wbd_imem_dat_o[21]
port 239 nsew signal output
rlabel metal2 s 83462 0 83518 800 6 wbd_imem_dat_o[22]
port 240 nsew signal output
rlabel metal2 s 84934 0 84990 800 6 wbd_imem_dat_o[23]
port 241 nsew signal output
rlabel metal2 s 86406 0 86462 800 6 wbd_imem_dat_o[24]
port 242 nsew signal output
rlabel metal2 s 87878 0 87934 800 6 wbd_imem_dat_o[25]
port 243 nsew signal output
rlabel metal2 s 89350 0 89406 800 6 wbd_imem_dat_o[26]
port 244 nsew signal output
rlabel metal2 s 90822 0 90878 800 6 wbd_imem_dat_o[27]
port 245 nsew signal output
rlabel metal2 s 92294 0 92350 800 6 wbd_imem_dat_o[28]
port 246 nsew signal output
rlabel metal2 s 93858 0 93914 800 6 wbd_imem_dat_o[29]
port 247 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 wbd_imem_dat_o[2]
port 248 nsew signal output
rlabel metal2 s 95330 0 95386 800 6 wbd_imem_dat_o[30]
port 249 nsew signal output
rlabel metal2 s 96802 0 96858 800 6 wbd_imem_dat_o[31]
port 250 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 wbd_imem_dat_o[3]
port 251 nsew signal output
rlabel metal2 s 56874 0 56930 800 6 wbd_imem_dat_o[4]
port 252 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 wbd_imem_dat_o[5]
port 253 nsew signal output
rlabel metal2 s 59818 0 59874 800 6 wbd_imem_dat_o[6]
port 254 nsew signal output
rlabel metal2 s 61290 0 61346 800 6 wbd_imem_dat_o[7]
port 255 nsew signal output
rlabel metal2 s 62762 0 62818 800 6 wbd_imem_dat_o[8]
port 256 nsew signal output
rlabel metal2 s 64234 0 64290 800 6 wbd_imem_dat_o[9]
port 257 nsew signal output
rlabel metal2 s 147034 0 147090 800 6 wbd_imem_err_i
port 258 nsew signal input
rlabel metal3 s 299200 233384 300000 233504 6 wbd_imem_sel_o[0]
port 259 nsew signal output
rlabel metal2 s 297730 0 297786 800 6 wbd_imem_sel_o[1]
port 260 nsew signal output
rlabel metal2 s 149978 239200 150034 240000 6 wbd_imem_sel_o[2]
port 261 nsew signal output
rlabel metal2 s 249982 239200 250038 240000 6 wbd_imem_sel_o[3]
port 262 nsew signal output
rlabel metal2 s 754 0 810 800 6 wbd_imem_stb_o
port 263 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 wbd_imem_we_o
port 264 nsew signal output
rlabel metal4 s 280688 2128 281008 237776 6 VPWR
port 265 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 237776 6 VPWR
port 266 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 237776 6 VPWR
port 267 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 237776 6 VPWR
port 268 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 237776 6 VPWR
port 269 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 237776 6 VPWR
port 270 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 237776 6 VPWR
port 271 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 237776 6 VPWR
port 272 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 237776 6 VPWR
port 273 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 237776 6 VPWR
port 274 nsew power bidirectional
rlabel metal5 s 1104 219750 298816 220070 6 VPWR
port 275 nsew power bidirectional
rlabel metal5 s 1104 189114 298816 189434 6 VPWR
port 276 nsew power bidirectional
rlabel metal5 s 1104 158478 298816 158798 6 VPWR
port 277 nsew power bidirectional
rlabel metal5 s 1104 127842 298816 128162 6 VPWR
port 278 nsew power bidirectional
rlabel metal5 s 1104 97206 298816 97526 6 VPWR
port 279 nsew power bidirectional
rlabel metal5 s 1104 66570 298816 66890 6 VPWR
port 280 nsew power bidirectional
rlabel metal5 s 1104 35934 298816 36254 6 VPWR
port 281 nsew power bidirectional
rlabel metal5 s 1104 5298 298816 5618 6 VPWR
port 282 nsew power bidirectional
rlabel metal4 s 296048 2128 296368 237776 6 VGND
port 283 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 237776 6 VGND
port 284 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 237776 6 VGND
port 285 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 237776 6 VGND
port 286 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 237776 6 VGND
port 287 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 237776 6 VGND
port 288 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 237776 6 VGND
port 289 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 237776 6 VGND
port 290 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 237776 6 VGND
port 291 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 237776 6 VGND
port 292 nsew ground bidirectional
rlabel metal5 s 1104 235068 298816 235388 6 VGND
port 293 nsew ground bidirectional
rlabel metal5 s 1104 204432 298816 204752 6 VGND
port 294 nsew ground bidirectional
rlabel metal5 s 1104 173796 298816 174116 6 VGND
port 295 nsew ground bidirectional
rlabel metal5 s 1104 143160 298816 143480 6 VGND
port 296 nsew ground bidirectional
rlabel metal5 s 1104 112524 298816 112844 6 VGND
port 297 nsew ground bidirectional
rlabel metal5 s 1104 81888 298816 82208 6 VGND
port 298 nsew ground bidirectional
rlabel metal5 s 1104 51252 298816 51572 6 VGND
port 299 nsew ground bidirectional
rlabel metal5 s 1104 20616 298816 20936 6 VGND
port 300 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 300000 240000
string LEFview TRUE
string GDS_FILE /project/openlane/syntacore/runs/syntacore/results/magic/scr1_top_wb.gds
string GDS_END 85558154
string GDS_START 301344
<< end >>

