magic
tech sky130A
magscale 1 2
timestamp 1623949457
<< obsli1 >>
rect 1380 1071 458620 19975
<< obsm1 >>
rect 658 8 459250 19984
<< metal2 >>
rect 662 19200 718 20000
rect 2042 19200 2098 20000
rect 3514 19200 3570 20000
rect 4986 19200 5042 20000
rect 6458 19200 6514 20000
rect 7930 19200 7986 20000
rect 9402 19200 9458 20000
rect 10874 19200 10930 20000
rect 12254 19200 12310 20000
rect 13726 19200 13782 20000
rect 15198 19200 15254 20000
rect 16670 19200 16726 20000
rect 18142 19200 18198 20000
rect 19614 19200 19670 20000
rect 21086 19200 21142 20000
rect 22558 19200 22614 20000
rect 23938 19200 23994 20000
rect 25410 19200 25466 20000
rect 26882 19200 26938 20000
rect 28354 19200 28410 20000
rect 29826 19200 29882 20000
rect 31298 19200 31354 20000
rect 32770 19200 32826 20000
rect 34242 19200 34298 20000
rect 35622 19200 35678 20000
rect 37094 19200 37150 20000
rect 38566 19200 38622 20000
rect 40038 19200 40094 20000
rect 41510 19200 41566 20000
rect 42982 19200 43038 20000
rect 44454 19200 44510 20000
rect 45926 19200 45982 20000
rect 47306 19200 47362 20000
rect 48778 19200 48834 20000
rect 50250 19200 50306 20000
rect 51722 19200 51778 20000
rect 53194 19200 53250 20000
rect 54666 19200 54722 20000
rect 56138 19200 56194 20000
rect 57610 19200 57666 20000
rect 58990 19200 59046 20000
rect 60462 19200 60518 20000
rect 61934 19200 61990 20000
rect 63406 19200 63462 20000
rect 64878 19200 64934 20000
rect 66350 19200 66406 20000
rect 67822 19200 67878 20000
rect 69294 19200 69350 20000
rect 70674 19200 70730 20000
rect 72146 19200 72202 20000
rect 73618 19200 73674 20000
rect 75090 19200 75146 20000
rect 76562 19200 76618 20000
rect 78034 19200 78090 20000
rect 79506 19200 79562 20000
rect 80978 19200 81034 20000
rect 82358 19200 82414 20000
rect 83830 19200 83886 20000
rect 85302 19200 85358 20000
rect 86774 19200 86830 20000
rect 88246 19200 88302 20000
rect 89718 19200 89774 20000
rect 91190 19200 91246 20000
rect 92662 19200 92718 20000
rect 94042 19200 94098 20000
rect 95514 19200 95570 20000
rect 96986 19200 97042 20000
rect 98458 19200 98514 20000
rect 99930 19200 99986 20000
rect 101402 19200 101458 20000
rect 102874 19200 102930 20000
rect 104254 19200 104310 20000
rect 105726 19200 105782 20000
rect 107198 19200 107254 20000
rect 108670 19200 108726 20000
rect 110142 19200 110198 20000
rect 111614 19200 111670 20000
rect 113086 19200 113142 20000
rect 114558 19200 114614 20000
rect 115938 19200 115994 20000
rect 117410 19200 117466 20000
rect 118882 19200 118938 20000
rect 120354 19200 120410 20000
rect 121826 19200 121882 20000
rect 123298 19200 123354 20000
rect 124770 19200 124826 20000
rect 126242 19200 126298 20000
rect 127622 19200 127678 20000
rect 129094 19200 129150 20000
rect 130566 19200 130622 20000
rect 132038 19200 132094 20000
rect 133510 19200 133566 20000
rect 134982 19200 135038 20000
rect 136454 19200 136510 20000
rect 137926 19200 137982 20000
rect 139306 19200 139362 20000
rect 140778 19200 140834 20000
rect 142250 19200 142306 20000
rect 143722 19200 143778 20000
rect 145194 19200 145250 20000
rect 146666 19200 146722 20000
rect 148138 19200 148194 20000
rect 149610 19200 149666 20000
rect 150990 19200 151046 20000
rect 152462 19200 152518 20000
rect 153934 19200 153990 20000
rect 155406 19200 155462 20000
rect 156878 19200 156934 20000
rect 158350 19200 158406 20000
rect 159822 19200 159878 20000
rect 161294 19200 161350 20000
rect 162674 19200 162730 20000
rect 164146 19200 164202 20000
rect 165618 19200 165674 20000
rect 167090 19200 167146 20000
rect 168562 19200 168618 20000
rect 170034 19200 170090 20000
rect 171506 19200 171562 20000
rect 172978 19200 173034 20000
rect 174358 19200 174414 20000
rect 175830 19200 175886 20000
rect 177302 19200 177358 20000
rect 178774 19200 178830 20000
rect 180246 19200 180302 20000
rect 181718 19200 181774 20000
rect 183190 19200 183246 20000
rect 184662 19200 184718 20000
rect 186042 19200 186098 20000
rect 187514 19200 187570 20000
rect 188986 19200 189042 20000
rect 190458 19200 190514 20000
rect 191930 19200 191986 20000
rect 193402 19200 193458 20000
rect 194874 19200 194930 20000
rect 196254 19200 196310 20000
rect 197726 19200 197782 20000
rect 199198 19200 199254 20000
rect 200670 19200 200726 20000
rect 202142 19200 202198 20000
rect 203614 19200 203670 20000
rect 205086 19200 205142 20000
rect 206558 19200 206614 20000
rect 207938 19200 207994 20000
rect 209410 19200 209466 20000
rect 210882 19200 210938 20000
rect 212354 19200 212410 20000
rect 213826 19200 213882 20000
rect 215298 19200 215354 20000
rect 216770 19200 216826 20000
rect 218242 19200 218298 20000
rect 219622 19200 219678 20000
rect 221094 19200 221150 20000
rect 222566 19200 222622 20000
rect 224038 19200 224094 20000
rect 225510 19200 225566 20000
rect 226982 19200 227038 20000
rect 228454 19200 228510 20000
rect 229926 19200 229982 20000
rect 231306 19200 231362 20000
rect 232778 19200 232834 20000
rect 234250 19200 234306 20000
rect 235722 19200 235778 20000
rect 237194 19200 237250 20000
rect 238666 19200 238722 20000
rect 240138 19200 240194 20000
rect 241610 19200 241666 20000
rect 242990 19200 243046 20000
rect 244462 19200 244518 20000
rect 245934 19200 245990 20000
rect 247406 19200 247462 20000
rect 248878 19200 248934 20000
rect 250350 19200 250406 20000
rect 251822 19200 251878 20000
rect 253294 19200 253350 20000
rect 254674 19200 254730 20000
rect 256146 19200 256202 20000
rect 257618 19200 257674 20000
rect 259090 19200 259146 20000
rect 260562 19200 260618 20000
rect 262034 19200 262090 20000
rect 263506 19200 263562 20000
rect 264978 19200 265034 20000
rect 266358 19200 266414 20000
rect 267830 19200 267886 20000
rect 269302 19200 269358 20000
rect 270774 19200 270830 20000
rect 272246 19200 272302 20000
rect 273718 19200 273774 20000
rect 275190 19200 275246 20000
rect 276662 19200 276718 20000
rect 278042 19200 278098 20000
rect 279514 19200 279570 20000
rect 280986 19200 281042 20000
rect 282458 19200 282514 20000
rect 283930 19200 283986 20000
rect 285402 19200 285458 20000
rect 286874 19200 286930 20000
rect 288254 19200 288310 20000
rect 289726 19200 289782 20000
rect 291198 19200 291254 20000
rect 292670 19200 292726 20000
rect 294142 19200 294198 20000
rect 295614 19200 295670 20000
rect 297086 19200 297142 20000
rect 298558 19200 298614 20000
rect 299938 19200 299994 20000
rect 301410 19200 301466 20000
rect 302882 19200 302938 20000
rect 304354 19200 304410 20000
rect 305826 19200 305882 20000
rect 307298 19200 307354 20000
rect 308770 19200 308826 20000
rect 310242 19200 310298 20000
rect 311622 19200 311678 20000
rect 313094 19200 313150 20000
rect 314566 19200 314622 20000
rect 316038 19200 316094 20000
rect 317510 19200 317566 20000
rect 318982 19200 319038 20000
rect 320454 19200 320510 20000
rect 321926 19200 321982 20000
rect 323306 19200 323362 20000
rect 324778 19200 324834 20000
rect 326250 19200 326306 20000
rect 327722 19200 327778 20000
rect 329194 19200 329250 20000
rect 330666 19200 330722 20000
rect 332138 19200 332194 20000
rect 333610 19200 333666 20000
rect 334990 19200 335046 20000
rect 336462 19200 336518 20000
rect 337934 19200 337990 20000
rect 339406 19200 339462 20000
rect 340878 19200 340934 20000
rect 342350 19200 342406 20000
rect 343822 19200 343878 20000
rect 345294 19200 345350 20000
rect 346674 19200 346730 20000
rect 348146 19200 348202 20000
rect 349618 19200 349674 20000
rect 351090 19200 351146 20000
rect 352562 19200 352618 20000
rect 354034 19200 354090 20000
rect 355506 19200 355562 20000
rect 356978 19200 357034 20000
rect 358358 19200 358414 20000
rect 359830 19200 359886 20000
rect 361302 19200 361358 20000
rect 362774 19200 362830 20000
rect 364246 19200 364302 20000
rect 365718 19200 365774 20000
rect 367190 19200 367246 20000
rect 368662 19200 368718 20000
rect 370042 19200 370098 20000
rect 371514 19200 371570 20000
rect 372986 19200 373042 20000
rect 374458 19200 374514 20000
rect 375930 19200 375986 20000
rect 377402 19200 377458 20000
rect 378874 19200 378930 20000
rect 380254 19200 380310 20000
rect 381726 19200 381782 20000
rect 383198 19200 383254 20000
rect 384670 19200 384726 20000
rect 386142 19200 386198 20000
rect 387614 19200 387670 20000
rect 389086 19200 389142 20000
rect 390558 19200 390614 20000
rect 391938 19200 391994 20000
rect 393410 19200 393466 20000
rect 394882 19200 394938 20000
rect 396354 19200 396410 20000
rect 397826 19200 397882 20000
rect 399298 19200 399354 20000
rect 400770 19200 400826 20000
rect 402242 19200 402298 20000
rect 403622 19200 403678 20000
rect 405094 19200 405150 20000
rect 406566 19200 406622 20000
rect 408038 19200 408094 20000
rect 409510 19200 409566 20000
rect 410982 19200 411038 20000
rect 412454 19200 412510 20000
rect 413926 19200 413982 20000
rect 415306 19200 415362 20000
rect 416778 19200 416834 20000
rect 418250 19200 418306 20000
rect 419722 19200 419778 20000
rect 421194 19200 421250 20000
rect 422666 19200 422722 20000
rect 424138 19200 424194 20000
rect 425610 19200 425666 20000
rect 426990 19200 427046 20000
rect 428462 19200 428518 20000
rect 429934 19200 429990 20000
rect 431406 19200 431462 20000
rect 432878 19200 432934 20000
rect 434350 19200 434406 20000
rect 435822 19200 435878 20000
rect 437294 19200 437350 20000
rect 438674 19200 438730 20000
rect 440146 19200 440202 20000
rect 441618 19200 441674 20000
rect 443090 19200 443146 20000
rect 444562 19200 444618 20000
rect 446034 19200 446090 20000
rect 447506 19200 447562 20000
rect 448978 19200 449034 20000
rect 450358 19200 450414 20000
rect 451830 19200 451886 20000
rect 453302 19200 453358 20000
rect 454774 19200 454830 20000
rect 456246 19200 456302 20000
rect 457718 19200 457774 20000
rect 459190 19200 459246 20000
rect 3350 1040 3410 18544
rect 11350 1040 11410 18544
rect 19350 1040 19410 18544
rect 27350 1040 27410 18544
rect 35350 1040 35410 18544
rect 43350 1040 43410 18544
rect 51350 1040 51410 18544
rect 59350 1040 59410 18544
rect 67350 1040 67410 18544
rect 75350 1040 75410 18544
rect 83350 1040 83410 18544
rect 91350 1040 91410 18544
rect 99350 1040 99410 18544
rect 107350 1040 107410 18544
rect 115350 1040 115410 18544
rect 123350 1040 123410 18544
rect 131350 1040 131410 18544
rect 139350 1040 139410 18544
rect 147350 1040 147410 18544
rect 155350 1040 155410 18544
rect 163350 1040 163410 18544
rect 171350 1040 171410 18544
rect 179350 1040 179410 18544
rect 187350 1040 187410 18544
rect 195350 1040 195410 18544
rect 203350 1040 203410 18544
rect 211350 1040 211410 18544
rect 219350 1040 219410 18544
rect 227350 1040 227410 18544
rect 235350 1040 235410 18544
rect 243350 1040 243410 18544
rect 251350 1040 251410 18544
rect 259350 1040 259410 18544
rect 267350 1040 267410 18544
rect 275350 1040 275410 18544
rect 283350 1040 283410 18544
rect 291350 1040 291410 18544
rect 299350 1040 299410 18544
rect 307350 1040 307410 18544
rect 315350 1040 315410 18544
rect 323350 1040 323410 18544
rect 331350 1040 331410 18544
rect 339350 1040 339410 18544
rect 347350 1040 347410 18544
rect 355350 1040 355410 18544
rect 363350 1040 363410 18544
rect 371350 1040 371410 18544
rect 379350 1040 379410 18544
rect 387350 1040 387410 18544
rect 395350 1040 395410 18544
rect 403350 1040 403410 18544
rect 411350 1040 411410 18544
rect 419350 1040 419410 18544
rect 427350 1040 427410 18544
rect 435350 1040 435410 18544
rect 443350 1040 443410 18544
rect 451350 1040 451410 18544
rect 662 0 718 800
rect 2042 0 2098 800
rect 3514 0 3570 800
rect 4986 0 5042 800
rect 6458 0 6514 800
rect 7930 0 7986 800
rect 9402 0 9458 800
rect 10874 0 10930 800
rect 12254 0 12310 800
rect 13726 0 13782 800
rect 15198 0 15254 800
rect 16670 0 16726 800
rect 18142 0 18198 800
rect 19614 0 19670 800
rect 21086 0 21142 800
rect 22558 0 22614 800
rect 23938 0 23994 800
rect 25410 0 25466 800
rect 26882 0 26938 800
rect 28354 0 28410 800
rect 29826 0 29882 800
rect 31298 0 31354 800
rect 32770 0 32826 800
rect 34242 0 34298 800
rect 35622 0 35678 800
rect 37094 0 37150 800
rect 38566 0 38622 800
rect 40038 0 40094 800
rect 41510 0 41566 800
rect 42982 0 43038 800
rect 44454 0 44510 800
rect 45926 0 45982 800
rect 47306 0 47362 800
rect 48778 0 48834 800
rect 50250 0 50306 800
rect 51722 0 51778 800
rect 53194 0 53250 800
rect 54666 0 54722 800
rect 56138 0 56194 800
rect 57610 0 57666 800
rect 58990 0 59046 800
rect 60462 0 60518 800
rect 61934 0 61990 800
rect 63406 0 63462 800
rect 64878 0 64934 800
rect 66350 0 66406 800
rect 67822 0 67878 800
rect 69294 0 69350 800
rect 70674 0 70730 800
rect 72146 0 72202 800
rect 73618 0 73674 800
rect 75090 0 75146 800
rect 76562 0 76618 800
rect 78034 0 78090 800
rect 79506 0 79562 800
rect 80978 0 81034 800
rect 82358 0 82414 800
rect 83830 0 83886 800
rect 85302 0 85358 800
rect 86774 0 86830 800
rect 88246 0 88302 800
rect 89718 0 89774 800
rect 91190 0 91246 800
rect 92662 0 92718 800
rect 94042 0 94098 800
rect 95514 0 95570 800
rect 96986 0 97042 800
rect 98458 0 98514 800
rect 99930 0 99986 800
rect 101402 0 101458 800
rect 102874 0 102930 800
rect 104254 0 104310 800
rect 105726 0 105782 800
rect 107198 0 107254 800
rect 108670 0 108726 800
rect 110142 0 110198 800
rect 111614 0 111670 800
rect 113086 0 113142 800
rect 114558 0 114614 800
rect 115938 0 115994 800
rect 117410 0 117466 800
rect 118882 0 118938 800
rect 120354 0 120410 800
rect 121826 0 121882 800
rect 123298 0 123354 800
rect 124770 0 124826 800
rect 126242 0 126298 800
rect 127622 0 127678 800
rect 129094 0 129150 800
rect 130566 0 130622 800
rect 132038 0 132094 800
rect 133510 0 133566 800
rect 134982 0 135038 800
rect 136454 0 136510 800
rect 137926 0 137982 800
rect 139306 0 139362 800
rect 140778 0 140834 800
rect 142250 0 142306 800
rect 143722 0 143778 800
rect 145194 0 145250 800
rect 146666 0 146722 800
rect 148138 0 148194 800
rect 149610 0 149666 800
rect 150990 0 151046 800
rect 152462 0 152518 800
rect 153934 0 153990 800
rect 155406 0 155462 800
rect 156878 0 156934 800
rect 158350 0 158406 800
rect 159822 0 159878 800
rect 161294 0 161350 800
rect 162674 0 162730 800
rect 164146 0 164202 800
rect 165618 0 165674 800
rect 167090 0 167146 800
rect 168562 0 168618 800
rect 170034 0 170090 800
rect 171506 0 171562 800
rect 172978 0 173034 800
rect 174358 0 174414 800
rect 175830 0 175886 800
rect 177302 0 177358 800
rect 178774 0 178830 800
rect 180246 0 180302 800
rect 181718 0 181774 800
rect 183190 0 183246 800
rect 184662 0 184718 800
rect 186042 0 186098 800
rect 187514 0 187570 800
rect 188986 0 189042 800
rect 190458 0 190514 800
rect 191930 0 191986 800
rect 193402 0 193458 800
rect 194874 0 194930 800
rect 196254 0 196310 800
rect 197726 0 197782 800
rect 199198 0 199254 800
rect 200670 0 200726 800
rect 202142 0 202198 800
rect 203614 0 203670 800
rect 205086 0 205142 800
rect 206558 0 206614 800
rect 207938 0 207994 800
rect 209410 0 209466 800
rect 210882 0 210938 800
rect 212354 0 212410 800
rect 213826 0 213882 800
rect 215298 0 215354 800
rect 216770 0 216826 800
rect 218242 0 218298 800
rect 219622 0 219678 800
rect 221094 0 221150 800
rect 222566 0 222622 800
rect 224038 0 224094 800
rect 225510 0 225566 800
rect 226982 0 227038 800
rect 228454 0 228510 800
rect 229926 0 229982 800
rect 231306 0 231362 800
rect 232778 0 232834 800
rect 234250 0 234306 800
rect 235722 0 235778 800
rect 237194 0 237250 800
rect 238666 0 238722 800
rect 240138 0 240194 800
rect 241610 0 241666 800
rect 242990 0 243046 800
rect 244462 0 244518 800
rect 245934 0 245990 800
rect 247406 0 247462 800
rect 248878 0 248934 800
rect 250350 0 250406 800
rect 251822 0 251878 800
rect 253294 0 253350 800
rect 254674 0 254730 800
rect 256146 0 256202 800
rect 257618 0 257674 800
rect 259090 0 259146 800
rect 260562 0 260618 800
rect 262034 0 262090 800
rect 263506 0 263562 800
rect 264978 0 265034 800
rect 266358 0 266414 800
rect 267830 0 267886 800
rect 269302 0 269358 800
rect 270774 0 270830 800
rect 272246 0 272302 800
rect 273718 0 273774 800
rect 275190 0 275246 800
rect 276662 0 276718 800
rect 278042 0 278098 800
rect 279514 0 279570 800
rect 280986 0 281042 800
rect 282458 0 282514 800
rect 283930 0 283986 800
rect 285402 0 285458 800
rect 286874 0 286930 800
rect 288254 0 288310 800
rect 289726 0 289782 800
rect 291198 0 291254 800
rect 292670 0 292726 800
rect 294142 0 294198 800
rect 295614 0 295670 800
rect 297086 0 297142 800
rect 298558 0 298614 800
rect 299938 0 299994 800
rect 301410 0 301466 800
rect 302882 0 302938 800
rect 304354 0 304410 800
rect 305826 0 305882 800
rect 307298 0 307354 800
rect 308770 0 308826 800
rect 310242 0 310298 800
rect 311622 0 311678 800
rect 313094 0 313150 800
rect 314566 0 314622 800
rect 316038 0 316094 800
rect 317510 0 317566 800
rect 318982 0 319038 800
rect 320454 0 320510 800
rect 321926 0 321982 800
rect 323306 0 323362 800
rect 324778 0 324834 800
rect 326250 0 326306 800
rect 327722 0 327778 800
rect 329194 0 329250 800
rect 330666 0 330722 800
rect 332138 0 332194 800
rect 333610 0 333666 800
rect 334990 0 335046 800
rect 336462 0 336518 800
rect 337934 0 337990 800
rect 339406 0 339462 800
rect 340878 0 340934 800
rect 342350 0 342406 800
rect 343822 0 343878 800
rect 345294 0 345350 800
rect 346674 0 346730 800
rect 348146 0 348202 800
rect 349618 0 349674 800
rect 351090 0 351146 800
rect 352562 0 352618 800
rect 354034 0 354090 800
rect 355506 0 355562 800
rect 356978 0 357034 800
rect 358358 0 358414 800
rect 359830 0 359886 800
rect 361302 0 361358 800
rect 362774 0 362830 800
rect 364246 0 364302 800
rect 365718 0 365774 800
rect 367190 0 367246 800
rect 368662 0 368718 800
rect 370042 0 370098 800
rect 371514 0 371570 800
rect 372986 0 373042 800
rect 374458 0 374514 800
rect 375930 0 375986 800
rect 377402 0 377458 800
rect 378874 0 378930 800
rect 380254 0 380310 800
rect 381726 0 381782 800
rect 383198 0 383254 800
rect 384670 0 384726 800
rect 386142 0 386198 800
rect 387614 0 387670 800
rect 389086 0 389142 800
rect 390558 0 390614 800
rect 391938 0 391994 800
rect 393410 0 393466 800
rect 394882 0 394938 800
rect 396354 0 396410 800
rect 397826 0 397882 800
rect 399298 0 399354 800
rect 400770 0 400826 800
rect 402242 0 402298 800
rect 403622 0 403678 800
rect 405094 0 405150 800
rect 406566 0 406622 800
rect 408038 0 408094 800
rect 409510 0 409566 800
rect 410982 0 411038 800
rect 412454 0 412510 800
rect 413926 0 413982 800
rect 415306 0 415362 800
rect 416778 0 416834 800
rect 418250 0 418306 800
rect 419722 0 419778 800
rect 421194 0 421250 800
rect 422666 0 422722 800
rect 424138 0 424194 800
rect 425610 0 425666 800
rect 426990 0 427046 800
rect 428462 0 428518 800
rect 429934 0 429990 800
rect 431406 0 431462 800
rect 432878 0 432934 800
rect 434350 0 434406 800
rect 435822 0 435878 800
rect 437294 0 437350 800
rect 438674 0 438730 800
rect 440146 0 440202 800
rect 441618 0 441674 800
rect 443090 0 443146 800
rect 444562 0 444618 800
rect 446034 0 446090 800
rect 447506 0 447562 800
rect 448978 0 449034 800
rect 450358 0 450414 800
rect 451830 0 451886 800
rect 453302 0 453358 800
rect 454774 0 454830 800
rect 456246 0 456302 800
rect 457718 0 457774 800
rect 459190 0 459246 800
<< obsm2 >>
rect 774 19144 1986 19990
rect 2154 19144 3458 19990
rect 3626 19144 4930 19990
rect 5098 19144 6402 19990
rect 6570 19144 7874 19990
rect 8042 19144 9346 19990
rect 9514 19144 10818 19990
rect 10986 19144 12198 19990
rect 12366 19144 13670 19990
rect 13838 19144 15142 19990
rect 15310 19144 16614 19990
rect 16782 19144 18086 19990
rect 18254 19144 19558 19990
rect 19726 19144 21030 19990
rect 21198 19144 22502 19990
rect 22670 19144 23882 19990
rect 24050 19144 25354 19990
rect 25522 19144 26826 19990
rect 26994 19144 28298 19990
rect 28466 19144 29770 19990
rect 29938 19144 31242 19990
rect 31410 19144 32714 19990
rect 32882 19144 34186 19990
rect 34354 19144 35566 19990
rect 35734 19144 37038 19990
rect 37206 19144 38510 19990
rect 38678 19144 39982 19990
rect 40150 19144 41454 19990
rect 41622 19144 42926 19990
rect 43094 19144 44398 19990
rect 44566 19144 45870 19990
rect 46038 19144 47250 19990
rect 47418 19144 48722 19990
rect 48890 19144 50194 19990
rect 50362 19144 51666 19990
rect 51834 19144 53138 19990
rect 53306 19144 54610 19990
rect 54778 19144 56082 19990
rect 56250 19144 57554 19990
rect 57722 19144 58934 19990
rect 59102 19144 60406 19990
rect 60574 19144 61878 19990
rect 62046 19144 63350 19990
rect 63518 19144 64822 19990
rect 64990 19144 66294 19990
rect 66462 19144 67766 19990
rect 67934 19144 69238 19990
rect 69406 19144 70618 19990
rect 70786 19144 72090 19990
rect 72258 19144 73562 19990
rect 73730 19144 75034 19990
rect 75202 19144 76506 19990
rect 76674 19144 77978 19990
rect 78146 19144 79450 19990
rect 79618 19144 80922 19990
rect 81090 19144 82302 19990
rect 82470 19144 83774 19990
rect 83942 19144 85246 19990
rect 85414 19144 86718 19990
rect 86886 19144 88190 19990
rect 88358 19144 89662 19990
rect 89830 19144 91134 19990
rect 91302 19144 92606 19990
rect 92774 19144 93986 19990
rect 94154 19144 95458 19990
rect 95626 19144 96930 19990
rect 97098 19144 98402 19990
rect 98570 19144 99874 19990
rect 100042 19144 101346 19990
rect 101514 19144 102818 19990
rect 102986 19144 104198 19990
rect 104366 19144 105670 19990
rect 105838 19144 107142 19990
rect 107310 19144 108614 19990
rect 108782 19144 110086 19990
rect 110254 19144 111558 19990
rect 111726 19144 113030 19990
rect 113198 19144 114502 19990
rect 114670 19144 115882 19990
rect 116050 19144 117354 19990
rect 117522 19144 118826 19990
rect 118994 19144 120298 19990
rect 120466 19144 121770 19990
rect 121938 19144 123242 19990
rect 123410 19144 124714 19990
rect 124882 19144 126186 19990
rect 126354 19144 127566 19990
rect 127734 19144 129038 19990
rect 129206 19144 130510 19990
rect 130678 19144 131982 19990
rect 132150 19144 133454 19990
rect 133622 19144 134926 19990
rect 135094 19144 136398 19990
rect 136566 19144 137870 19990
rect 138038 19144 139250 19990
rect 139418 19144 140722 19990
rect 140890 19144 142194 19990
rect 142362 19144 143666 19990
rect 143834 19144 145138 19990
rect 145306 19144 146610 19990
rect 146778 19144 148082 19990
rect 148250 19144 149554 19990
rect 149722 19144 150934 19990
rect 151102 19144 152406 19990
rect 152574 19144 153878 19990
rect 154046 19144 155350 19990
rect 155518 19144 156822 19990
rect 156990 19144 158294 19990
rect 158462 19144 159766 19990
rect 159934 19144 161238 19990
rect 161406 19144 162618 19990
rect 162786 19144 164090 19990
rect 164258 19144 165562 19990
rect 165730 19144 167034 19990
rect 167202 19144 168506 19990
rect 168674 19144 169978 19990
rect 170146 19144 171450 19990
rect 171618 19144 172922 19990
rect 173090 19144 174302 19990
rect 174470 19144 175774 19990
rect 175942 19144 177246 19990
rect 177414 19144 178718 19990
rect 178886 19144 180190 19990
rect 180358 19144 181662 19990
rect 181830 19144 183134 19990
rect 183302 19144 184606 19990
rect 184774 19144 185986 19990
rect 186154 19144 187458 19990
rect 187626 19144 188930 19990
rect 189098 19144 190402 19990
rect 190570 19144 191874 19990
rect 192042 19144 193346 19990
rect 193514 19144 194818 19990
rect 194986 19144 196198 19990
rect 196366 19144 197670 19990
rect 197838 19144 199142 19990
rect 199310 19144 200614 19990
rect 200782 19144 202086 19990
rect 202254 19144 203558 19990
rect 203726 19144 205030 19990
rect 205198 19144 206502 19990
rect 206670 19144 207882 19990
rect 208050 19144 209354 19990
rect 209522 19144 210826 19990
rect 210994 19144 212298 19990
rect 212466 19144 213770 19990
rect 213938 19144 215242 19990
rect 215410 19144 216714 19990
rect 216882 19144 218186 19990
rect 218354 19144 219566 19990
rect 219734 19144 221038 19990
rect 221206 19144 222510 19990
rect 222678 19144 223982 19990
rect 224150 19144 225454 19990
rect 225622 19144 226926 19990
rect 227094 19144 228398 19990
rect 228566 19144 229870 19990
rect 230038 19144 231250 19990
rect 231418 19144 232722 19990
rect 232890 19144 234194 19990
rect 234362 19144 235666 19990
rect 235834 19144 237138 19990
rect 237306 19144 238610 19990
rect 238778 19144 240082 19990
rect 240250 19144 241554 19990
rect 241722 19144 242934 19990
rect 243102 19144 244406 19990
rect 244574 19144 245878 19990
rect 246046 19144 247350 19990
rect 247518 19144 248822 19990
rect 248990 19144 250294 19990
rect 250462 19144 251766 19990
rect 251934 19144 253238 19990
rect 253406 19144 254618 19990
rect 254786 19144 256090 19990
rect 256258 19144 257562 19990
rect 257730 19144 259034 19990
rect 259202 19144 260506 19990
rect 260674 19144 261978 19990
rect 262146 19144 263450 19990
rect 263618 19144 264922 19990
rect 265090 19144 266302 19990
rect 266470 19144 267774 19990
rect 267942 19144 269246 19990
rect 269414 19144 270718 19990
rect 270886 19144 272190 19990
rect 272358 19144 273662 19990
rect 273830 19144 275134 19990
rect 275302 19144 276606 19990
rect 276774 19144 277986 19990
rect 278154 19144 279458 19990
rect 279626 19144 280930 19990
rect 281098 19144 282402 19990
rect 282570 19144 283874 19990
rect 284042 19144 285346 19990
rect 285514 19144 286818 19990
rect 286986 19144 288198 19990
rect 288366 19144 289670 19990
rect 289838 19144 291142 19990
rect 291310 19144 292614 19990
rect 292782 19144 294086 19990
rect 294254 19144 295558 19990
rect 295726 19144 297030 19990
rect 297198 19144 298502 19990
rect 298670 19144 299882 19990
rect 300050 19144 301354 19990
rect 301522 19144 302826 19990
rect 302994 19144 304298 19990
rect 304466 19144 305770 19990
rect 305938 19144 307242 19990
rect 307410 19144 308714 19990
rect 308882 19144 310186 19990
rect 310354 19144 311566 19990
rect 311734 19144 313038 19990
rect 313206 19144 314510 19990
rect 314678 19144 315982 19990
rect 316150 19144 317454 19990
rect 317622 19144 318926 19990
rect 319094 19144 320398 19990
rect 320566 19144 321870 19990
rect 322038 19144 323250 19990
rect 323418 19144 324722 19990
rect 324890 19144 326194 19990
rect 326362 19144 327666 19990
rect 327834 19144 329138 19990
rect 329306 19144 330610 19990
rect 330778 19144 332082 19990
rect 332250 19144 333554 19990
rect 333722 19144 334934 19990
rect 335102 19144 336406 19990
rect 336574 19144 337878 19990
rect 338046 19144 339350 19990
rect 339518 19144 340822 19990
rect 340990 19144 342294 19990
rect 342462 19144 343766 19990
rect 343934 19144 345238 19990
rect 345406 19144 346618 19990
rect 346786 19144 348090 19990
rect 348258 19144 349562 19990
rect 349730 19144 351034 19990
rect 351202 19144 352506 19990
rect 352674 19144 353978 19990
rect 354146 19144 355450 19990
rect 355618 19144 356922 19990
rect 357090 19144 358302 19990
rect 358470 19144 359774 19990
rect 359942 19144 361246 19990
rect 361414 19144 362718 19990
rect 362886 19144 364190 19990
rect 364358 19144 365662 19990
rect 365830 19144 367134 19990
rect 367302 19144 368606 19990
rect 368774 19144 369986 19990
rect 370154 19144 371458 19990
rect 371626 19144 372930 19990
rect 373098 19144 374402 19990
rect 374570 19144 375874 19990
rect 376042 19144 377346 19990
rect 377514 19144 378818 19990
rect 378986 19144 380198 19990
rect 380366 19144 381670 19990
rect 381838 19144 383142 19990
rect 383310 19144 384614 19990
rect 384782 19144 386086 19990
rect 386254 19144 387558 19990
rect 387726 19144 389030 19990
rect 389198 19144 390502 19990
rect 390670 19144 391882 19990
rect 392050 19144 393354 19990
rect 393522 19144 394826 19990
rect 394994 19144 396298 19990
rect 396466 19144 397770 19990
rect 397938 19144 399242 19990
rect 399410 19144 400714 19990
rect 400882 19144 402186 19990
rect 402354 19144 403566 19990
rect 403734 19144 405038 19990
rect 405206 19144 406510 19990
rect 406678 19144 407982 19990
rect 408150 19144 409454 19990
rect 409622 19144 410926 19990
rect 411094 19144 412398 19990
rect 412566 19144 413870 19990
rect 414038 19144 415250 19990
rect 415418 19144 416722 19990
rect 416890 19144 418194 19990
rect 418362 19144 419666 19990
rect 419834 19144 421138 19990
rect 421306 19144 422610 19990
rect 422778 19144 424082 19990
rect 424250 19144 425554 19990
rect 425722 19144 426934 19990
rect 427102 19144 428406 19990
rect 428574 19144 429878 19990
rect 430046 19144 431350 19990
rect 431518 19144 432822 19990
rect 432990 19144 434294 19990
rect 434462 19144 435766 19990
rect 435934 19144 437238 19990
rect 437406 19144 438618 19990
rect 438786 19144 440090 19990
rect 440258 19144 441562 19990
rect 441730 19144 443034 19990
rect 443202 19144 444506 19990
rect 444674 19144 445978 19990
rect 446146 19144 447450 19990
rect 447618 19144 448922 19990
rect 449090 19144 450302 19990
rect 450470 19144 451774 19990
rect 451942 19144 453246 19990
rect 453414 19144 454718 19990
rect 454886 19144 456190 19990
rect 456358 19144 457662 19990
rect 457830 19144 459134 19990
rect 664 18600 459246 19144
rect 664 984 3294 18600
rect 3466 984 11294 18600
rect 11466 984 19294 18600
rect 19466 984 27294 18600
rect 27466 984 35294 18600
rect 35466 984 43294 18600
rect 43466 984 51294 18600
rect 51466 984 59294 18600
rect 59466 984 67294 18600
rect 67466 984 75294 18600
rect 75466 984 83294 18600
rect 83466 984 91294 18600
rect 91466 984 99294 18600
rect 99466 984 107294 18600
rect 107466 984 115294 18600
rect 115466 984 123294 18600
rect 123466 984 131294 18600
rect 131466 984 139294 18600
rect 139466 984 147294 18600
rect 147466 984 155294 18600
rect 155466 984 163294 18600
rect 163466 984 171294 18600
rect 171466 984 179294 18600
rect 179466 984 187294 18600
rect 187466 984 195294 18600
rect 195466 984 203294 18600
rect 203466 984 211294 18600
rect 211466 984 219294 18600
rect 219466 984 227294 18600
rect 227466 984 235294 18600
rect 235466 984 243294 18600
rect 243466 984 251294 18600
rect 251466 984 259294 18600
rect 259466 984 267294 18600
rect 267466 984 275294 18600
rect 275466 984 283294 18600
rect 283466 984 291294 18600
rect 291466 984 299294 18600
rect 299466 984 307294 18600
rect 307466 984 315294 18600
rect 315466 984 323294 18600
rect 323466 984 331294 18600
rect 331466 984 339294 18600
rect 339466 984 347294 18600
rect 347466 984 355294 18600
rect 355466 984 363294 18600
rect 363466 984 371294 18600
rect 371466 984 379294 18600
rect 379466 984 387294 18600
rect 387466 984 395294 18600
rect 395466 984 403294 18600
rect 403466 984 411294 18600
rect 411466 984 419294 18600
rect 419466 984 427294 18600
rect 427466 984 435294 18600
rect 435466 984 443294 18600
rect 443466 984 451294 18600
rect 451466 984 459246 18600
rect 664 856 459246 984
rect 774 2 1986 856
rect 2154 2 3458 856
rect 3626 2 4930 856
rect 5098 2 6402 856
rect 6570 2 7874 856
rect 8042 2 9346 856
rect 9514 2 10818 856
rect 10986 2 12198 856
rect 12366 2 13670 856
rect 13838 2 15142 856
rect 15310 2 16614 856
rect 16782 2 18086 856
rect 18254 2 19558 856
rect 19726 2 21030 856
rect 21198 2 22502 856
rect 22670 2 23882 856
rect 24050 2 25354 856
rect 25522 2 26826 856
rect 26994 2 28298 856
rect 28466 2 29770 856
rect 29938 2 31242 856
rect 31410 2 32714 856
rect 32882 2 34186 856
rect 34354 2 35566 856
rect 35734 2 37038 856
rect 37206 2 38510 856
rect 38678 2 39982 856
rect 40150 2 41454 856
rect 41622 2 42926 856
rect 43094 2 44398 856
rect 44566 2 45870 856
rect 46038 2 47250 856
rect 47418 2 48722 856
rect 48890 2 50194 856
rect 50362 2 51666 856
rect 51834 2 53138 856
rect 53306 2 54610 856
rect 54778 2 56082 856
rect 56250 2 57554 856
rect 57722 2 58934 856
rect 59102 2 60406 856
rect 60574 2 61878 856
rect 62046 2 63350 856
rect 63518 2 64822 856
rect 64990 2 66294 856
rect 66462 2 67766 856
rect 67934 2 69238 856
rect 69406 2 70618 856
rect 70786 2 72090 856
rect 72258 2 73562 856
rect 73730 2 75034 856
rect 75202 2 76506 856
rect 76674 2 77978 856
rect 78146 2 79450 856
rect 79618 2 80922 856
rect 81090 2 82302 856
rect 82470 2 83774 856
rect 83942 2 85246 856
rect 85414 2 86718 856
rect 86886 2 88190 856
rect 88358 2 89662 856
rect 89830 2 91134 856
rect 91302 2 92606 856
rect 92774 2 93986 856
rect 94154 2 95458 856
rect 95626 2 96930 856
rect 97098 2 98402 856
rect 98570 2 99874 856
rect 100042 2 101346 856
rect 101514 2 102818 856
rect 102986 2 104198 856
rect 104366 2 105670 856
rect 105838 2 107142 856
rect 107310 2 108614 856
rect 108782 2 110086 856
rect 110254 2 111558 856
rect 111726 2 113030 856
rect 113198 2 114502 856
rect 114670 2 115882 856
rect 116050 2 117354 856
rect 117522 2 118826 856
rect 118994 2 120298 856
rect 120466 2 121770 856
rect 121938 2 123242 856
rect 123410 2 124714 856
rect 124882 2 126186 856
rect 126354 2 127566 856
rect 127734 2 129038 856
rect 129206 2 130510 856
rect 130678 2 131982 856
rect 132150 2 133454 856
rect 133622 2 134926 856
rect 135094 2 136398 856
rect 136566 2 137870 856
rect 138038 2 139250 856
rect 139418 2 140722 856
rect 140890 2 142194 856
rect 142362 2 143666 856
rect 143834 2 145138 856
rect 145306 2 146610 856
rect 146778 2 148082 856
rect 148250 2 149554 856
rect 149722 2 150934 856
rect 151102 2 152406 856
rect 152574 2 153878 856
rect 154046 2 155350 856
rect 155518 2 156822 856
rect 156990 2 158294 856
rect 158462 2 159766 856
rect 159934 2 161238 856
rect 161406 2 162618 856
rect 162786 2 164090 856
rect 164258 2 165562 856
rect 165730 2 167034 856
rect 167202 2 168506 856
rect 168674 2 169978 856
rect 170146 2 171450 856
rect 171618 2 172922 856
rect 173090 2 174302 856
rect 174470 2 175774 856
rect 175942 2 177246 856
rect 177414 2 178718 856
rect 178886 2 180190 856
rect 180358 2 181662 856
rect 181830 2 183134 856
rect 183302 2 184606 856
rect 184774 2 185986 856
rect 186154 2 187458 856
rect 187626 2 188930 856
rect 189098 2 190402 856
rect 190570 2 191874 856
rect 192042 2 193346 856
rect 193514 2 194818 856
rect 194986 2 196198 856
rect 196366 2 197670 856
rect 197838 2 199142 856
rect 199310 2 200614 856
rect 200782 2 202086 856
rect 202254 2 203558 856
rect 203726 2 205030 856
rect 205198 2 206502 856
rect 206670 2 207882 856
rect 208050 2 209354 856
rect 209522 2 210826 856
rect 210994 2 212298 856
rect 212466 2 213770 856
rect 213938 2 215242 856
rect 215410 2 216714 856
rect 216882 2 218186 856
rect 218354 2 219566 856
rect 219734 2 221038 856
rect 221206 2 222510 856
rect 222678 2 223982 856
rect 224150 2 225454 856
rect 225622 2 226926 856
rect 227094 2 228398 856
rect 228566 2 229870 856
rect 230038 2 231250 856
rect 231418 2 232722 856
rect 232890 2 234194 856
rect 234362 2 235666 856
rect 235834 2 237138 856
rect 237306 2 238610 856
rect 238778 2 240082 856
rect 240250 2 241554 856
rect 241722 2 242934 856
rect 243102 2 244406 856
rect 244574 2 245878 856
rect 246046 2 247350 856
rect 247518 2 248822 856
rect 248990 2 250294 856
rect 250462 2 251766 856
rect 251934 2 253238 856
rect 253406 2 254618 856
rect 254786 2 256090 856
rect 256258 2 257562 856
rect 257730 2 259034 856
rect 259202 2 260506 856
rect 260674 2 261978 856
rect 262146 2 263450 856
rect 263618 2 264922 856
rect 265090 2 266302 856
rect 266470 2 267774 856
rect 267942 2 269246 856
rect 269414 2 270718 856
rect 270886 2 272190 856
rect 272358 2 273662 856
rect 273830 2 275134 856
rect 275302 2 276606 856
rect 276774 2 277986 856
rect 278154 2 279458 856
rect 279626 2 280930 856
rect 281098 2 282402 856
rect 282570 2 283874 856
rect 284042 2 285346 856
rect 285514 2 286818 856
rect 286986 2 288198 856
rect 288366 2 289670 856
rect 289838 2 291142 856
rect 291310 2 292614 856
rect 292782 2 294086 856
rect 294254 2 295558 856
rect 295726 2 297030 856
rect 297198 2 298502 856
rect 298670 2 299882 856
rect 300050 2 301354 856
rect 301522 2 302826 856
rect 302994 2 304298 856
rect 304466 2 305770 856
rect 305938 2 307242 856
rect 307410 2 308714 856
rect 308882 2 310186 856
rect 310354 2 311566 856
rect 311734 2 313038 856
rect 313206 2 314510 856
rect 314678 2 315982 856
rect 316150 2 317454 856
rect 317622 2 318926 856
rect 319094 2 320398 856
rect 320566 2 321870 856
rect 322038 2 323250 856
rect 323418 2 324722 856
rect 324890 2 326194 856
rect 326362 2 327666 856
rect 327834 2 329138 856
rect 329306 2 330610 856
rect 330778 2 332082 856
rect 332250 2 333554 856
rect 333722 2 334934 856
rect 335102 2 336406 856
rect 336574 2 337878 856
rect 338046 2 339350 856
rect 339518 2 340822 856
rect 340990 2 342294 856
rect 342462 2 343766 856
rect 343934 2 345238 856
rect 345406 2 346618 856
rect 346786 2 348090 856
rect 348258 2 349562 856
rect 349730 2 351034 856
rect 351202 2 352506 856
rect 352674 2 353978 856
rect 354146 2 355450 856
rect 355618 2 356922 856
rect 357090 2 358302 856
rect 358470 2 359774 856
rect 359942 2 361246 856
rect 361414 2 362718 856
rect 362886 2 364190 856
rect 364358 2 365662 856
rect 365830 2 367134 856
rect 367302 2 368606 856
rect 368774 2 369986 856
rect 370154 2 371458 856
rect 371626 2 372930 856
rect 373098 2 374402 856
rect 374570 2 375874 856
rect 376042 2 377346 856
rect 377514 2 378818 856
rect 378986 2 380198 856
rect 380366 2 381670 856
rect 381838 2 383142 856
rect 383310 2 384614 856
rect 384782 2 386086 856
rect 386254 2 387558 856
rect 387726 2 389030 856
rect 389198 2 390502 856
rect 390670 2 391882 856
rect 392050 2 393354 856
rect 393522 2 394826 856
rect 394994 2 396298 856
rect 396466 2 397770 856
rect 397938 2 399242 856
rect 399410 2 400714 856
rect 400882 2 402186 856
rect 402354 2 403566 856
rect 403734 2 405038 856
rect 405206 2 406510 856
rect 406678 2 407982 856
rect 408150 2 409454 856
rect 409622 2 410926 856
rect 411094 2 412398 856
rect 412566 2 413870 856
rect 414038 2 415250 856
rect 415418 2 416722 856
rect 416890 2 418194 856
rect 418362 2 419666 856
rect 419834 2 421138 856
rect 421306 2 422610 856
rect 422778 2 424082 856
rect 424250 2 425554 856
rect 425722 2 426934 856
rect 427102 2 428406 856
rect 428574 2 429878 856
rect 430046 2 431350 856
rect 431518 2 432822 856
rect 432990 2 434294 856
rect 434462 2 435766 856
rect 435934 2 437238 856
rect 437406 2 438618 856
rect 438786 2 440090 856
rect 440258 2 441562 856
rect 441730 2 443034 856
rect 443202 2 444506 856
rect 444674 2 445978 856
rect 446146 2 447450 856
rect 447618 2 448922 856
rect 449090 2 450302 856
rect 450470 2 451774 856
rect 451942 2 453246 856
rect 453414 2 454718 856
rect 454886 2 456190 856
rect 456358 2 457662 856
rect 457830 2 459134 856
<< metal3 >>
rect 1380 17410 458620 17470
rect 1380 16330 458620 16390
rect 1380 15250 458620 15310
rect 459200 14832 460000 14952
rect 1380 14170 458620 14230
rect 1380 13090 458620 13150
rect 1380 12010 458620 12070
rect 1380 10930 458620 10990
rect 1380 9850 458620 9910
rect 1380 8770 458620 8830
rect 1380 7690 458620 7750
rect 1380 6610 458620 6670
rect 1380 5530 458620 5590
rect 459200 4904 460000 5024
rect 1380 4450 458620 4510
rect 1380 3370 458620 3430
rect 1380 2290 458620 2350
rect 1380 1210 458620 1270
<< obsm3 >>
rect 3347 17550 459251 19957
rect 458700 17330 459251 17550
rect 3347 16470 459251 17330
rect 458700 16250 459251 16470
rect 3347 15390 459251 16250
rect 458700 15170 459251 15390
rect 3347 15032 459251 15170
rect 3347 14752 459120 15032
rect 3347 14310 459251 14752
rect 458700 14090 459251 14310
rect 3347 13230 459251 14090
rect 458700 13010 459251 13230
rect 3347 12150 459251 13010
rect 458700 11930 459251 12150
rect 3347 11070 459251 11930
rect 458700 10850 459251 11070
rect 3347 9990 459251 10850
rect 458700 9770 459251 9990
rect 3347 8910 459251 9770
rect 458700 8690 459251 8910
rect 3347 7830 459251 8690
rect 458700 7610 459251 7830
rect 3347 6750 459251 7610
rect 458700 6530 459251 6750
rect 3347 5670 459251 6530
rect 458700 5450 459251 5670
rect 3347 5104 459251 5450
rect 3347 4824 459120 5104
rect 3347 4590 459251 4824
rect 458700 4370 459251 4590
rect 3347 3510 459251 4370
rect 458700 3290 459251 3510
rect 3347 2430 459251 3290
rect 458700 2210 459251 2430
rect 3347 1350 459251 2210
rect 458700 1130 459251 1350
rect 3347 35 459251 1130
<< labels >>
rlabel metal3 s 459200 4904 460000 5024 6 clk_i
port 1 nsew signal input
rlabel metal2 s 149610 19200 149666 20000 6 m0_wbd_ack_o
port 2 nsew signal output
rlabel metal2 s 3514 19200 3570 20000 6 m0_wbd_adr_i[0]
port 3 nsew signal input
rlabel metal2 s 18142 19200 18198 20000 6 m0_wbd_adr_i[10]
port 4 nsew signal input
rlabel metal2 s 19614 19200 19670 20000 6 m0_wbd_adr_i[11]
port 5 nsew signal input
rlabel metal2 s 21086 19200 21142 20000 6 m0_wbd_adr_i[12]
port 6 nsew signal input
rlabel metal2 s 22558 19200 22614 20000 6 m0_wbd_adr_i[13]
port 7 nsew signal input
rlabel metal2 s 23938 19200 23994 20000 6 m0_wbd_adr_i[14]
port 8 nsew signal input
rlabel metal2 s 25410 19200 25466 20000 6 m0_wbd_adr_i[15]
port 9 nsew signal input
rlabel metal2 s 26882 19200 26938 20000 6 m0_wbd_adr_i[16]
port 10 nsew signal input
rlabel metal2 s 28354 19200 28410 20000 6 m0_wbd_adr_i[17]
port 11 nsew signal input
rlabel metal2 s 29826 19200 29882 20000 6 m0_wbd_adr_i[18]
port 12 nsew signal input
rlabel metal2 s 31298 19200 31354 20000 6 m0_wbd_adr_i[19]
port 13 nsew signal input
rlabel metal2 s 4986 19200 5042 20000 6 m0_wbd_adr_i[1]
port 14 nsew signal input
rlabel metal2 s 32770 19200 32826 20000 6 m0_wbd_adr_i[20]
port 15 nsew signal input
rlabel metal2 s 34242 19200 34298 20000 6 m0_wbd_adr_i[21]
port 16 nsew signal input
rlabel metal2 s 35622 19200 35678 20000 6 m0_wbd_adr_i[22]
port 17 nsew signal input
rlabel metal2 s 37094 19200 37150 20000 6 m0_wbd_adr_i[23]
port 18 nsew signal input
rlabel metal2 s 38566 19200 38622 20000 6 m0_wbd_adr_i[24]
port 19 nsew signal input
rlabel metal2 s 40038 19200 40094 20000 6 m0_wbd_adr_i[25]
port 20 nsew signal input
rlabel metal2 s 41510 19200 41566 20000 6 m0_wbd_adr_i[26]
port 21 nsew signal input
rlabel metal2 s 42982 19200 43038 20000 6 m0_wbd_adr_i[27]
port 22 nsew signal input
rlabel metal2 s 44454 19200 44510 20000 6 m0_wbd_adr_i[28]
port 23 nsew signal input
rlabel metal2 s 45926 19200 45982 20000 6 m0_wbd_adr_i[29]
port 24 nsew signal input
rlabel metal2 s 6458 19200 6514 20000 6 m0_wbd_adr_i[2]
port 25 nsew signal input
rlabel metal2 s 47306 19200 47362 20000 6 m0_wbd_adr_i[30]
port 26 nsew signal input
rlabel metal2 s 48778 19200 48834 20000 6 m0_wbd_adr_i[31]
port 27 nsew signal input
rlabel metal2 s 7930 19200 7986 20000 6 m0_wbd_adr_i[3]
port 28 nsew signal input
rlabel metal2 s 9402 19200 9458 20000 6 m0_wbd_adr_i[4]
port 29 nsew signal input
rlabel metal2 s 10874 19200 10930 20000 6 m0_wbd_adr_i[5]
port 30 nsew signal input
rlabel metal2 s 12254 19200 12310 20000 6 m0_wbd_adr_i[6]
port 31 nsew signal input
rlabel metal2 s 13726 19200 13782 20000 6 m0_wbd_adr_i[7]
port 32 nsew signal input
rlabel metal2 s 15198 19200 15254 20000 6 m0_wbd_adr_i[8]
port 33 nsew signal input
rlabel metal2 s 16670 19200 16726 20000 6 m0_wbd_adr_i[9]
port 34 nsew signal input
rlabel metal2 s 152462 19200 152518 20000 6 m0_wbd_cyc_i
port 35 nsew signal input
rlabel metal2 s 56138 19200 56194 20000 6 m0_wbd_dat_i[0]
port 36 nsew signal input
rlabel metal2 s 70674 19200 70730 20000 6 m0_wbd_dat_i[10]
port 37 nsew signal input
rlabel metal2 s 72146 19200 72202 20000 6 m0_wbd_dat_i[11]
port 38 nsew signal input
rlabel metal2 s 73618 19200 73674 20000 6 m0_wbd_dat_i[12]
port 39 nsew signal input
rlabel metal2 s 75090 19200 75146 20000 6 m0_wbd_dat_i[13]
port 40 nsew signal input
rlabel metal2 s 76562 19200 76618 20000 6 m0_wbd_dat_i[14]
port 41 nsew signal input
rlabel metal2 s 78034 19200 78090 20000 6 m0_wbd_dat_i[15]
port 42 nsew signal input
rlabel metal2 s 79506 19200 79562 20000 6 m0_wbd_dat_i[16]
port 43 nsew signal input
rlabel metal2 s 80978 19200 81034 20000 6 m0_wbd_dat_i[17]
port 44 nsew signal input
rlabel metal2 s 82358 19200 82414 20000 6 m0_wbd_dat_i[18]
port 45 nsew signal input
rlabel metal2 s 83830 19200 83886 20000 6 m0_wbd_dat_i[19]
port 46 nsew signal input
rlabel metal2 s 57610 19200 57666 20000 6 m0_wbd_dat_i[1]
port 47 nsew signal input
rlabel metal2 s 85302 19200 85358 20000 6 m0_wbd_dat_i[20]
port 48 nsew signal input
rlabel metal2 s 86774 19200 86830 20000 6 m0_wbd_dat_i[21]
port 49 nsew signal input
rlabel metal2 s 88246 19200 88302 20000 6 m0_wbd_dat_i[22]
port 50 nsew signal input
rlabel metal2 s 89718 19200 89774 20000 6 m0_wbd_dat_i[23]
port 51 nsew signal input
rlabel metal2 s 91190 19200 91246 20000 6 m0_wbd_dat_i[24]
port 52 nsew signal input
rlabel metal2 s 92662 19200 92718 20000 6 m0_wbd_dat_i[25]
port 53 nsew signal input
rlabel metal2 s 94042 19200 94098 20000 6 m0_wbd_dat_i[26]
port 54 nsew signal input
rlabel metal2 s 95514 19200 95570 20000 6 m0_wbd_dat_i[27]
port 55 nsew signal input
rlabel metal2 s 96986 19200 97042 20000 6 m0_wbd_dat_i[28]
port 56 nsew signal input
rlabel metal2 s 98458 19200 98514 20000 6 m0_wbd_dat_i[29]
port 57 nsew signal input
rlabel metal2 s 58990 19200 59046 20000 6 m0_wbd_dat_i[2]
port 58 nsew signal input
rlabel metal2 s 99930 19200 99986 20000 6 m0_wbd_dat_i[30]
port 59 nsew signal input
rlabel metal2 s 101402 19200 101458 20000 6 m0_wbd_dat_i[31]
port 60 nsew signal input
rlabel metal2 s 60462 19200 60518 20000 6 m0_wbd_dat_i[3]
port 61 nsew signal input
rlabel metal2 s 61934 19200 61990 20000 6 m0_wbd_dat_i[4]
port 62 nsew signal input
rlabel metal2 s 63406 19200 63462 20000 6 m0_wbd_dat_i[5]
port 63 nsew signal input
rlabel metal2 s 64878 19200 64934 20000 6 m0_wbd_dat_i[6]
port 64 nsew signal input
rlabel metal2 s 66350 19200 66406 20000 6 m0_wbd_dat_i[7]
port 65 nsew signal input
rlabel metal2 s 67822 19200 67878 20000 6 m0_wbd_dat_i[8]
port 66 nsew signal input
rlabel metal2 s 69294 19200 69350 20000 6 m0_wbd_dat_i[9]
port 67 nsew signal input
rlabel metal2 s 102874 19200 102930 20000 6 m0_wbd_dat_o[0]
port 68 nsew signal output
rlabel metal2 s 117410 19200 117466 20000 6 m0_wbd_dat_o[10]
port 69 nsew signal output
rlabel metal2 s 118882 19200 118938 20000 6 m0_wbd_dat_o[11]
port 70 nsew signal output
rlabel metal2 s 120354 19200 120410 20000 6 m0_wbd_dat_o[12]
port 71 nsew signal output
rlabel metal2 s 121826 19200 121882 20000 6 m0_wbd_dat_o[13]
port 72 nsew signal output
rlabel metal2 s 123298 19200 123354 20000 6 m0_wbd_dat_o[14]
port 73 nsew signal output
rlabel metal2 s 124770 19200 124826 20000 6 m0_wbd_dat_o[15]
port 74 nsew signal output
rlabel metal2 s 126242 19200 126298 20000 6 m0_wbd_dat_o[16]
port 75 nsew signal output
rlabel metal2 s 127622 19200 127678 20000 6 m0_wbd_dat_o[17]
port 76 nsew signal output
rlabel metal2 s 129094 19200 129150 20000 6 m0_wbd_dat_o[18]
port 77 nsew signal output
rlabel metal2 s 130566 19200 130622 20000 6 m0_wbd_dat_o[19]
port 78 nsew signal output
rlabel metal2 s 104254 19200 104310 20000 6 m0_wbd_dat_o[1]
port 79 nsew signal output
rlabel metal2 s 132038 19200 132094 20000 6 m0_wbd_dat_o[20]
port 80 nsew signal output
rlabel metal2 s 133510 19200 133566 20000 6 m0_wbd_dat_o[21]
port 81 nsew signal output
rlabel metal2 s 134982 19200 135038 20000 6 m0_wbd_dat_o[22]
port 82 nsew signal output
rlabel metal2 s 136454 19200 136510 20000 6 m0_wbd_dat_o[23]
port 83 nsew signal output
rlabel metal2 s 137926 19200 137982 20000 6 m0_wbd_dat_o[24]
port 84 nsew signal output
rlabel metal2 s 139306 19200 139362 20000 6 m0_wbd_dat_o[25]
port 85 nsew signal output
rlabel metal2 s 140778 19200 140834 20000 6 m0_wbd_dat_o[26]
port 86 nsew signal output
rlabel metal2 s 142250 19200 142306 20000 6 m0_wbd_dat_o[27]
port 87 nsew signal output
rlabel metal2 s 143722 19200 143778 20000 6 m0_wbd_dat_o[28]
port 88 nsew signal output
rlabel metal2 s 145194 19200 145250 20000 6 m0_wbd_dat_o[29]
port 89 nsew signal output
rlabel metal2 s 105726 19200 105782 20000 6 m0_wbd_dat_o[2]
port 90 nsew signal output
rlabel metal2 s 146666 19200 146722 20000 6 m0_wbd_dat_o[30]
port 91 nsew signal output
rlabel metal2 s 148138 19200 148194 20000 6 m0_wbd_dat_o[31]
port 92 nsew signal output
rlabel metal2 s 107198 19200 107254 20000 6 m0_wbd_dat_o[3]
port 93 nsew signal output
rlabel metal2 s 108670 19200 108726 20000 6 m0_wbd_dat_o[4]
port 94 nsew signal output
rlabel metal2 s 110142 19200 110198 20000 6 m0_wbd_dat_o[5]
port 95 nsew signal output
rlabel metal2 s 111614 19200 111670 20000 6 m0_wbd_dat_o[6]
port 96 nsew signal output
rlabel metal2 s 113086 19200 113142 20000 6 m0_wbd_dat_o[7]
port 97 nsew signal output
rlabel metal2 s 114558 19200 114614 20000 6 m0_wbd_dat_o[8]
port 98 nsew signal output
rlabel metal2 s 115938 19200 115994 20000 6 m0_wbd_dat_o[9]
port 99 nsew signal output
rlabel metal2 s 150990 19200 151046 20000 6 m0_wbd_err_o
port 100 nsew signal output
rlabel metal2 s 50250 19200 50306 20000 6 m0_wbd_sel_i[0]
port 101 nsew signal input
rlabel metal2 s 51722 19200 51778 20000 6 m0_wbd_sel_i[1]
port 102 nsew signal input
rlabel metal2 s 53194 19200 53250 20000 6 m0_wbd_sel_i[2]
port 103 nsew signal input
rlabel metal2 s 54666 19200 54722 20000 6 m0_wbd_sel_i[3]
port 104 nsew signal input
rlabel metal2 s 662 19200 718 20000 6 m0_wbd_stb_i
port 105 nsew signal input
rlabel metal2 s 2042 19200 2098 20000 6 m0_wbd_we_i
port 106 nsew signal input
rlabel metal2 s 302882 19200 302938 20000 6 m1_wbd_ack_o
port 107 nsew signal output
rlabel metal2 s 156878 19200 156934 20000 6 m1_wbd_adr_i[0]
port 108 nsew signal input
rlabel metal2 s 171506 19200 171562 20000 6 m1_wbd_adr_i[10]
port 109 nsew signal input
rlabel metal2 s 172978 19200 173034 20000 6 m1_wbd_adr_i[11]
port 110 nsew signal input
rlabel metal2 s 174358 19200 174414 20000 6 m1_wbd_adr_i[12]
port 111 nsew signal input
rlabel metal2 s 175830 19200 175886 20000 6 m1_wbd_adr_i[13]
port 112 nsew signal input
rlabel metal2 s 177302 19200 177358 20000 6 m1_wbd_adr_i[14]
port 113 nsew signal input
rlabel metal2 s 178774 19200 178830 20000 6 m1_wbd_adr_i[15]
port 114 nsew signal input
rlabel metal2 s 180246 19200 180302 20000 6 m1_wbd_adr_i[16]
port 115 nsew signal input
rlabel metal2 s 181718 19200 181774 20000 6 m1_wbd_adr_i[17]
port 116 nsew signal input
rlabel metal2 s 183190 19200 183246 20000 6 m1_wbd_adr_i[18]
port 117 nsew signal input
rlabel metal2 s 184662 19200 184718 20000 6 m1_wbd_adr_i[19]
port 118 nsew signal input
rlabel metal2 s 158350 19200 158406 20000 6 m1_wbd_adr_i[1]
port 119 nsew signal input
rlabel metal2 s 186042 19200 186098 20000 6 m1_wbd_adr_i[20]
port 120 nsew signal input
rlabel metal2 s 187514 19200 187570 20000 6 m1_wbd_adr_i[21]
port 121 nsew signal input
rlabel metal2 s 188986 19200 189042 20000 6 m1_wbd_adr_i[22]
port 122 nsew signal input
rlabel metal2 s 190458 19200 190514 20000 6 m1_wbd_adr_i[23]
port 123 nsew signal input
rlabel metal2 s 191930 19200 191986 20000 6 m1_wbd_adr_i[24]
port 124 nsew signal input
rlabel metal2 s 193402 19200 193458 20000 6 m1_wbd_adr_i[25]
port 125 nsew signal input
rlabel metal2 s 194874 19200 194930 20000 6 m1_wbd_adr_i[26]
port 126 nsew signal input
rlabel metal2 s 196254 19200 196310 20000 6 m1_wbd_adr_i[27]
port 127 nsew signal input
rlabel metal2 s 197726 19200 197782 20000 6 m1_wbd_adr_i[28]
port 128 nsew signal input
rlabel metal2 s 199198 19200 199254 20000 6 m1_wbd_adr_i[29]
port 129 nsew signal input
rlabel metal2 s 159822 19200 159878 20000 6 m1_wbd_adr_i[2]
port 130 nsew signal input
rlabel metal2 s 200670 19200 200726 20000 6 m1_wbd_adr_i[30]
port 131 nsew signal input
rlabel metal2 s 202142 19200 202198 20000 6 m1_wbd_adr_i[31]
port 132 nsew signal input
rlabel metal2 s 161294 19200 161350 20000 6 m1_wbd_adr_i[3]
port 133 nsew signal input
rlabel metal2 s 162674 19200 162730 20000 6 m1_wbd_adr_i[4]
port 134 nsew signal input
rlabel metal2 s 164146 19200 164202 20000 6 m1_wbd_adr_i[5]
port 135 nsew signal input
rlabel metal2 s 165618 19200 165674 20000 6 m1_wbd_adr_i[6]
port 136 nsew signal input
rlabel metal2 s 167090 19200 167146 20000 6 m1_wbd_adr_i[7]
port 137 nsew signal input
rlabel metal2 s 168562 19200 168618 20000 6 m1_wbd_adr_i[8]
port 138 nsew signal input
rlabel metal2 s 170034 19200 170090 20000 6 m1_wbd_adr_i[9]
port 139 nsew signal input
rlabel metal2 s 305826 19200 305882 20000 6 m1_wbd_cyc_i
port 140 nsew signal input
rlabel metal2 s 209410 19200 209466 20000 6 m1_wbd_dat_i[0]
port 141 nsew signal input
rlabel metal2 s 224038 19200 224094 20000 6 m1_wbd_dat_i[10]
port 142 nsew signal input
rlabel metal2 s 225510 19200 225566 20000 6 m1_wbd_dat_i[11]
port 143 nsew signal input
rlabel metal2 s 226982 19200 227038 20000 6 m1_wbd_dat_i[12]
port 144 nsew signal input
rlabel metal2 s 228454 19200 228510 20000 6 m1_wbd_dat_i[13]
port 145 nsew signal input
rlabel metal2 s 229926 19200 229982 20000 6 m1_wbd_dat_i[14]
port 146 nsew signal input
rlabel metal2 s 231306 19200 231362 20000 6 m1_wbd_dat_i[15]
port 147 nsew signal input
rlabel metal2 s 232778 19200 232834 20000 6 m1_wbd_dat_i[16]
port 148 nsew signal input
rlabel metal2 s 234250 19200 234306 20000 6 m1_wbd_dat_i[17]
port 149 nsew signal input
rlabel metal2 s 235722 19200 235778 20000 6 m1_wbd_dat_i[18]
port 150 nsew signal input
rlabel metal2 s 237194 19200 237250 20000 6 m1_wbd_dat_i[19]
port 151 nsew signal input
rlabel metal2 s 210882 19200 210938 20000 6 m1_wbd_dat_i[1]
port 152 nsew signal input
rlabel metal2 s 238666 19200 238722 20000 6 m1_wbd_dat_i[20]
port 153 nsew signal input
rlabel metal2 s 240138 19200 240194 20000 6 m1_wbd_dat_i[21]
port 154 nsew signal input
rlabel metal2 s 241610 19200 241666 20000 6 m1_wbd_dat_i[22]
port 155 nsew signal input
rlabel metal2 s 242990 19200 243046 20000 6 m1_wbd_dat_i[23]
port 156 nsew signal input
rlabel metal2 s 244462 19200 244518 20000 6 m1_wbd_dat_i[24]
port 157 nsew signal input
rlabel metal2 s 245934 19200 245990 20000 6 m1_wbd_dat_i[25]
port 158 nsew signal input
rlabel metal2 s 247406 19200 247462 20000 6 m1_wbd_dat_i[26]
port 159 nsew signal input
rlabel metal2 s 248878 19200 248934 20000 6 m1_wbd_dat_i[27]
port 160 nsew signal input
rlabel metal2 s 250350 19200 250406 20000 6 m1_wbd_dat_i[28]
port 161 nsew signal input
rlabel metal2 s 251822 19200 251878 20000 6 m1_wbd_dat_i[29]
port 162 nsew signal input
rlabel metal2 s 212354 19200 212410 20000 6 m1_wbd_dat_i[2]
port 163 nsew signal input
rlabel metal2 s 253294 19200 253350 20000 6 m1_wbd_dat_i[30]
port 164 nsew signal input
rlabel metal2 s 254674 19200 254730 20000 6 m1_wbd_dat_i[31]
port 165 nsew signal input
rlabel metal2 s 213826 19200 213882 20000 6 m1_wbd_dat_i[3]
port 166 nsew signal input
rlabel metal2 s 215298 19200 215354 20000 6 m1_wbd_dat_i[4]
port 167 nsew signal input
rlabel metal2 s 216770 19200 216826 20000 6 m1_wbd_dat_i[5]
port 168 nsew signal input
rlabel metal2 s 218242 19200 218298 20000 6 m1_wbd_dat_i[6]
port 169 nsew signal input
rlabel metal2 s 219622 19200 219678 20000 6 m1_wbd_dat_i[7]
port 170 nsew signal input
rlabel metal2 s 221094 19200 221150 20000 6 m1_wbd_dat_i[8]
port 171 nsew signal input
rlabel metal2 s 222566 19200 222622 20000 6 m1_wbd_dat_i[9]
port 172 nsew signal input
rlabel metal2 s 256146 19200 256202 20000 6 m1_wbd_dat_o[0]
port 173 nsew signal output
rlabel metal2 s 270774 19200 270830 20000 6 m1_wbd_dat_o[10]
port 174 nsew signal output
rlabel metal2 s 272246 19200 272302 20000 6 m1_wbd_dat_o[11]
port 175 nsew signal output
rlabel metal2 s 273718 19200 273774 20000 6 m1_wbd_dat_o[12]
port 176 nsew signal output
rlabel metal2 s 275190 19200 275246 20000 6 m1_wbd_dat_o[13]
port 177 nsew signal output
rlabel metal2 s 276662 19200 276718 20000 6 m1_wbd_dat_o[14]
port 178 nsew signal output
rlabel metal2 s 278042 19200 278098 20000 6 m1_wbd_dat_o[15]
port 179 nsew signal output
rlabel metal2 s 279514 19200 279570 20000 6 m1_wbd_dat_o[16]
port 180 nsew signal output
rlabel metal2 s 280986 19200 281042 20000 6 m1_wbd_dat_o[17]
port 181 nsew signal output
rlabel metal2 s 282458 19200 282514 20000 6 m1_wbd_dat_o[18]
port 182 nsew signal output
rlabel metal2 s 283930 19200 283986 20000 6 m1_wbd_dat_o[19]
port 183 nsew signal output
rlabel metal2 s 257618 19200 257674 20000 6 m1_wbd_dat_o[1]
port 184 nsew signal output
rlabel metal2 s 285402 19200 285458 20000 6 m1_wbd_dat_o[20]
port 185 nsew signal output
rlabel metal2 s 286874 19200 286930 20000 6 m1_wbd_dat_o[21]
port 186 nsew signal output
rlabel metal2 s 288254 19200 288310 20000 6 m1_wbd_dat_o[22]
port 187 nsew signal output
rlabel metal2 s 289726 19200 289782 20000 6 m1_wbd_dat_o[23]
port 188 nsew signal output
rlabel metal2 s 291198 19200 291254 20000 6 m1_wbd_dat_o[24]
port 189 nsew signal output
rlabel metal2 s 292670 19200 292726 20000 6 m1_wbd_dat_o[25]
port 190 nsew signal output
rlabel metal2 s 294142 19200 294198 20000 6 m1_wbd_dat_o[26]
port 191 nsew signal output
rlabel metal2 s 295614 19200 295670 20000 6 m1_wbd_dat_o[27]
port 192 nsew signal output
rlabel metal2 s 297086 19200 297142 20000 6 m1_wbd_dat_o[28]
port 193 nsew signal output
rlabel metal2 s 298558 19200 298614 20000 6 m1_wbd_dat_o[29]
port 194 nsew signal output
rlabel metal2 s 259090 19200 259146 20000 6 m1_wbd_dat_o[2]
port 195 nsew signal output
rlabel metal2 s 299938 19200 299994 20000 6 m1_wbd_dat_o[30]
port 196 nsew signal output
rlabel metal2 s 301410 19200 301466 20000 6 m1_wbd_dat_o[31]
port 197 nsew signal output
rlabel metal2 s 260562 19200 260618 20000 6 m1_wbd_dat_o[3]
port 198 nsew signal output
rlabel metal2 s 262034 19200 262090 20000 6 m1_wbd_dat_o[4]
port 199 nsew signal output
rlabel metal2 s 263506 19200 263562 20000 6 m1_wbd_dat_o[5]
port 200 nsew signal output
rlabel metal2 s 264978 19200 265034 20000 6 m1_wbd_dat_o[6]
port 201 nsew signal output
rlabel metal2 s 266358 19200 266414 20000 6 m1_wbd_dat_o[7]
port 202 nsew signal output
rlabel metal2 s 267830 19200 267886 20000 6 m1_wbd_dat_o[8]
port 203 nsew signal output
rlabel metal2 s 269302 19200 269358 20000 6 m1_wbd_dat_o[9]
port 204 nsew signal output
rlabel metal2 s 304354 19200 304410 20000 6 m1_wbd_err_o
port 205 nsew signal output
rlabel metal2 s 203614 19200 203670 20000 6 m1_wbd_sel_i[0]
port 206 nsew signal input
rlabel metal2 s 205086 19200 205142 20000 6 m1_wbd_sel_i[1]
port 207 nsew signal input
rlabel metal2 s 206558 19200 206614 20000 6 m1_wbd_sel_i[2]
port 208 nsew signal input
rlabel metal2 s 207938 19200 207994 20000 6 m1_wbd_sel_i[3]
port 209 nsew signal input
rlabel metal2 s 153934 19200 153990 20000 6 m1_wbd_stb_i
port 210 nsew signal input
rlabel metal2 s 155406 19200 155462 20000 6 m1_wbd_we_i
port 211 nsew signal input
rlabel metal2 s 456246 19200 456302 20000 6 m2_wbd_ack_o
port 212 nsew signal output
rlabel metal2 s 310242 19200 310298 20000 6 m2_wbd_adr_i[0]
port 213 nsew signal input
rlabel metal2 s 324778 19200 324834 20000 6 m2_wbd_adr_i[10]
port 214 nsew signal input
rlabel metal2 s 326250 19200 326306 20000 6 m2_wbd_adr_i[11]
port 215 nsew signal input
rlabel metal2 s 327722 19200 327778 20000 6 m2_wbd_adr_i[12]
port 216 nsew signal input
rlabel metal2 s 329194 19200 329250 20000 6 m2_wbd_adr_i[13]
port 217 nsew signal input
rlabel metal2 s 330666 19200 330722 20000 6 m2_wbd_adr_i[14]
port 218 nsew signal input
rlabel metal2 s 332138 19200 332194 20000 6 m2_wbd_adr_i[15]
port 219 nsew signal input
rlabel metal2 s 333610 19200 333666 20000 6 m2_wbd_adr_i[16]
port 220 nsew signal input
rlabel metal2 s 334990 19200 335046 20000 6 m2_wbd_adr_i[17]
port 221 nsew signal input
rlabel metal2 s 336462 19200 336518 20000 6 m2_wbd_adr_i[18]
port 222 nsew signal input
rlabel metal2 s 337934 19200 337990 20000 6 m2_wbd_adr_i[19]
port 223 nsew signal input
rlabel metal2 s 311622 19200 311678 20000 6 m2_wbd_adr_i[1]
port 224 nsew signal input
rlabel metal2 s 339406 19200 339462 20000 6 m2_wbd_adr_i[20]
port 225 nsew signal input
rlabel metal2 s 340878 19200 340934 20000 6 m2_wbd_adr_i[21]
port 226 nsew signal input
rlabel metal2 s 342350 19200 342406 20000 6 m2_wbd_adr_i[22]
port 227 nsew signal input
rlabel metal2 s 343822 19200 343878 20000 6 m2_wbd_adr_i[23]
port 228 nsew signal input
rlabel metal2 s 345294 19200 345350 20000 6 m2_wbd_adr_i[24]
port 229 nsew signal input
rlabel metal2 s 346674 19200 346730 20000 6 m2_wbd_adr_i[25]
port 230 nsew signal input
rlabel metal2 s 348146 19200 348202 20000 6 m2_wbd_adr_i[26]
port 231 nsew signal input
rlabel metal2 s 349618 19200 349674 20000 6 m2_wbd_adr_i[27]
port 232 nsew signal input
rlabel metal2 s 351090 19200 351146 20000 6 m2_wbd_adr_i[28]
port 233 nsew signal input
rlabel metal2 s 352562 19200 352618 20000 6 m2_wbd_adr_i[29]
port 234 nsew signal input
rlabel metal2 s 313094 19200 313150 20000 6 m2_wbd_adr_i[2]
port 235 nsew signal input
rlabel metal2 s 354034 19200 354090 20000 6 m2_wbd_adr_i[30]
port 236 nsew signal input
rlabel metal2 s 355506 19200 355562 20000 6 m2_wbd_adr_i[31]
port 237 nsew signal input
rlabel metal2 s 314566 19200 314622 20000 6 m2_wbd_adr_i[3]
port 238 nsew signal input
rlabel metal2 s 316038 19200 316094 20000 6 m2_wbd_adr_i[4]
port 239 nsew signal input
rlabel metal2 s 317510 19200 317566 20000 6 m2_wbd_adr_i[5]
port 240 nsew signal input
rlabel metal2 s 318982 19200 319038 20000 6 m2_wbd_adr_i[6]
port 241 nsew signal input
rlabel metal2 s 320454 19200 320510 20000 6 m2_wbd_adr_i[7]
port 242 nsew signal input
rlabel metal2 s 321926 19200 321982 20000 6 m2_wbd_adr_i[8]
port 243 nsew signal input
rlabel metal2 s 323306 19200 323362 20000 6 m2_wbd_adr_i[9]
port 244 nsew signal input
rlabel metal2 s 459190 19200 459246 20000 6 m2_wbd_cyc_i
port 245 nsew signal input
rlabel metal2 s 362774 19200 362830 20000 6 m2_wbd_dat_i[0]
port 246 nsew signal input
rlabel metal2 s 377402 19200 377458 20000 6 m2_wbd_dat_i[10]
port 247 nsew signal input
rlabel metal2 s 378874 19200 378930 20000 6 m2_wbd_dat_i[11]
port 248 nsew signal input
rlabel metal2 s 380254 19200 380310 20000 6 m2_wbd_dat_i[12]
port 249 nsew signal input
rlabel metal2 s 381726 19200 381782 20000 6 m2_wbd_dat_i[13]
port 250 nsew signal input
rlabel metal2 s 383198 19200 383254 20000 6 m2_wbd_dat_i[14]
port 251 nsew signal input
rlabel metal2 s 384670 19200 384726 20000 6 m2_wbd_dat_i[15]
port 252 nsew signal input
rlabel metal2 s 386142 19200 386198 20000 6 m2_wbd_dat_i[16]
port 253 nsew signal input
rlabel metal2 s 387614 19200 387670 20000 6 m2_wbd_dat_i[17]
port 254 nsew signal input
rlabel metal2 s 389086 19200 389142 20000 6 m2_wbd_dat_i[18]
port 255 nsew signal input
rlabel metal2 s 390558 19200 390614 20000 6 m2_wbd_dat_i[19]
port 256 nsew signal input
rlabel metal2 s 364246 19200 364302 20000 6 m2_wbd_dat_i[1]
port 257 nsew signal input
rlabel metal2 s 391938 19200 391994 20000 6 m2_wbd_dat_i[20]
port 258 nsew signal input
rlabel metal2 s 393410 19200 393466 20000 6 m2_wbd_dat_i[21]
port 259 nsew signal input
rlabel metal2 s 394882 19200 394938 20000 6 m2_wbd_dat_i[22]
port 260 nsew signal input
rlabel metal2 s 396354 19200 396410 20000 6 m2_wbd_dat_i[23]
port 261 nsew signal input
rlabel metal2 s 397826 19200 397882 20000 6 m2_wbd_dat_i[24]
port 262 nsew signal input
rlabel metal2 s 399298 19200 399354 20000 6 m2_wbd_dat_i[25]
port 263 nsew signal input
rlabel metal2 s 400770 19200 400826 20000 6 m2_wbd_dat_i[26]
port 264 nsew signal input
rlabel metal2 s 402242 19200 402298 20000 6 m2_wbd_dat_i[27]
port 265 nsew signal input
rlabel metal2 s 403622 19200 403678 20000 6 m2_wbd_dat_i[28]
port 266 nsew signal input
rlabel metal2 s 405094 19200 405150 20000 6 m2_wbd_dat_i[29]
port 267 nsew signal input
rlabel metal2 s 365718 19200 365774 20000 6 m2_wbd_dat_i[2]
port 268 nsew signal input
rlabel metal2 s 406566 19200 406622 20000 6 m2_wbd_dat_i[30]
port 269 nsew signal input
rlabel metal2 s 408038 19200 408094 20000 6 m2_wbd_dat_i[31]
port 270 nsew signal input
rlabel metal2 s 367190 19200 367246 20000 6 m2_wbd_dat_i[3]
port 271 nsew signal input
rlabel metal2 s 368662 19200 368718 20000 6 m2_wbd_dat_i[4]
port 272 nsew signal input
rlabel metal2 s 370042 19200 370098 20000 6 m2_wbd_dat_i[5]
port 273 nsew signal input
rlabel metal2 s 371514 19200 371570 20000 6 m2_wbd_dat_i[6]
port 274 nsew signal input
rlabel metal2 s 372986 19200 373042 20000 6 m2_wbd_dat_i[7]
port 275 nsew signal input
rlabel metal2 s 374458 19200 374514 20000 6 m2_wbd_dat_i[8]
port 276 nsew signal input
rlabel metal2 s 375930 19200 375986 20000 6 m2_wbd_dat_i[9]
port 277 nsew signal input
rlabel metal2 s 409510 19200 409566 20000 6 m2_wbd_dat_o[0]
port 278 nsew signal output
rlabel metal2 s 424138 19200 424194 20000 6 m2_wbd_dat_o[10]
port 279 nsew signal output
rlabel metal2 s 425610 19200 425666 20000 6 m2_wbd_dat_o[11]
port 280 nsew signal output
rlabel metal2 s 426990 19200 427046 20000 6 m2_wbd_dat_o[12]
port 281 nsew signal output
rlabel metal2 s 428462 19200 428518 20000 6 m2_wbd_dat_o[13]
port 282 nsew signal output
rlabel metal2 s 429934 19200 429990 20000 6 m2_wbd_dat_o[14]
port 283 nsew signal output
rlabel metal2 s 431406 19200 431462 20000 6 m2_wbd_dat_o[15]
port 284 nsew signal output
rlabel metal2 s 432878 19200 432934 20000 6 m2_wbd_dat_o[16]
port 285 nsew signal output
rlabel metal2 s 434350 19200 434406 20000 6 m2_wbd_dat_o[17]
port 286 nsew signal output
rlabel metal2 s 435822 19200 435878 20000 6 m2_wbd_dat_o[18]
port 287 nsew signal output
rlabel metal2 s 437294 19200 437350 20000 6 m2_wbd_dat_o[19]
port 288 nsew signal output
rlabel metal2 s 410982 19200 411038 20000 6 m2_wbd_dat_o[1]
port 289 nsew signal output
rlabel metal2 s 438674 19200 438730 20000 6 m2_wbd_dat_o[20]
port 290 nsew signal output
rlabel metal2 s 440146 19200 440202 20000 6 m2_wbd_dat_o[21]
port 291 nsew signal output
rlabel metal2 s 441618 19200 441674 20000 6 m2_wbd_dat_o[22]
port 292 nsew signal output
rlabel metal2 s 443090 19200 443146 20000 6 m2_wbd_dat_o[23]
port 293 nsew signal output
rlabel metal2 s 444562 19200 444618 20000 6 m2_wbd_dat_o[24]
port 294 nsew signal output
rlabel metal2 s 446034 19200 446090 20000 6 m2_wbd_dat_o[25]
port 295 nsew signal output
rlabel metal2 s 447506 19200 447562 20000 6 m2_wbd_dat_o[26]
port 296 nsew signal output
rlabel metal2 s 448978 19200 449034 20000 6 m2_wbd_dat_o[27]
port 297 nsew signal output
rlabel metal2 s 450358 19200 450414 20000 6 m2_wbd_dat_o[28]
port 298 nsew signal output
rlabel metal2 s 451830 19200 451886 20000 6 m2_wbd_dat_o[29]
port 299 nsew signal output
rlabel metal2 s 412454 19200 412510 20000 6 m2_wbd_dat_o[2]
port 300 nsew signal output
rlabel metal2 s 453302 19200 453358 20000 6 m2_wbd_dat_o[30]
port 301 nsew signal output
rlabel metal2 s 454774 19200 454830 20000 6 m2_wbd_dat_o[31]
port 302 nsew signal output
rlabel metal2 s 413926 19200 413982 20000 6 m2_wbd_dat_o[3]
port 303 nsew signal output
rlabel metal2 s 415306 19200 415362 20000 6 m2_wbd_dat_o[4]
port 304 nsew signal output
rlabel metal2 s 416778 19200 416834 20000 6 m2_wbd_dat_o[5]
port 305 nsew signal output
rlabel metal2 s 418250 19200 418306 20000 6 m2_wbd_dat_o[6]
port 306 nsew signal output
rlabel metal2 s 419722 19200 419778 20000 6 m2_wbd_dat_o[7]
port 307 nsew signal output
rlabel metal2 s 421194 19200 421250 20000 6 m2_wbd_dat_o[8]
port 308 nsew signal output
rlabel metal2 s 422666 19200 422722 20000 6 m2_wbd_dat_o[9]
port 309 nsew signal output
rlabel metal2 s 457718 19200 457774 20000 6 m2_wbd_err_o
port 310 nsew signal output
rlabel metal2 s 356978 19200 357034 20000 6 m2_wbd_sel_i[0]
port 311 nsew signal input
rlabel metal2 s 358358 19200 358414 20000 6 m2_wbd_sel_i[1]
port 312 nsew signal input
rlabel metal2 s 359830 19200 359886 20000 6 m2_wbd_sel_i[2]
port 313 nsew signal input
rlabel metal2 s 361302 19200 361358 20000 6 m2_wbd_sel_i[3]
port 314 nsew signal input
rlabel metal2 s 307298 19200 307354 20000 6 m2_wbd_stb_i
port 315 nsew signal input
rlabel metal2 s 308770 19200 308826 20000 6 m2_wbd_we_i
port 316 nsew signal input
rlabel metal3 s 459200 14832 460000 14952 6 rst_n
port 317 nsew signal input
rlabel metal2 s 149610 0 149666 800 6 s0_wbd_ack_i
port 318 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 s0_wbd_adr_o[0]
port 319 nsew signal output
rlabel metal2 s 18142 0 18198 800 6 s0_wbd_adr_o[10]
port 320 nsew signal output
rlabel metal2 s 19614 0 19670 800 6 s0_wbd_adr_o[11]
port 321 nsew signal output
rlabel metal2 s 21086 0 21142 800 6 s0_wbd_adr_o[12]
port 322 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 s0_wbd_adr_o[13]
port 323 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 s0_wbd_adr_o[14]
port 324 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 s0_wbd_adr_o[15]
port 325 nsew signal output
rlabel metal2 s 26882 0 26938 800 6 s0_wbd_adr_o[16]
port 326 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 s0_wbd_adr_o[17]
port 327 nsew signal output
rlabel metal2 s 29826 0 29882 800 6 s0_wbd_adr_o[18]
port 328 nsew signal output
rlabel metal2 s 31298 0 31354 800 6 s0_wbd_adr_o[19]
port 329 nsew signal output
rlabel metal2 s 4986 0 5042 800 6 s0_wbd_adr_o[1]
port 330 nsew signal output
rlabel metal2 s 32770 0 32826 800 6 s0_wbd_adr_o[20]
port 331 nsew signal output
rlabel metal2 s 34242 0 34298 800 6 s0_wbd_adr_o[21]
port 332 nsew signal output
rlabel metal2 s 35622 0 35678 800 6 s0_wbd_adr_o[22]
port 333 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 s0_wbd_adr_o[23]
port 334 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 s0_wbd_adr_o[24]
port 335 nsew signal output
rlabel metal2 s 40038 0 40094 800 6 s0_wbd_adr_o[25]
port 336 nsew signal output
rlabel metal2 s 41510 0 41566 800 6 s0_wbd_adr_o[26]
port 337 nsew signal output
rlabel metal2 s 42982 0 43038 800 6 s0_wbd_adr_o[27]
port 338 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 s0_wbd_adr_o[28]
port 339 nsew signal output
rlabel metal2 s 45926 0 45982 800 6 s0_wbd_adr_o[29]
port 340 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 s0_wbd_adr_o[2]
port 341 nsew signal output
rlabel metal2 s 47306 0 47362 800 6 s0_wbd_adr_o[30]
port 342 nsew signal output
rlabel metal2 s 48778 0 48834 800 6 s0_wbd_adr_o[31]
port 343 nsew signal output
rlabel metal2 s 7930 0 7986 800 6 s0_wbd_adr_o[3]
port 344 nsew signal output
rlabel metal2 s 9402 0 9458 800 6 s0_wbd_adr_o[4]
port 345 nsew signal output
rlabel metal2 s 10874 0 10930 800 6 s0_wbd_adr_o[5]
port 346 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 s0_wbd_adr_o[6]
port 347 nsew signal output
rlabel metal2 s 13726 0 13782 800 6 s0_wbd_adr_o[7]
port 348 nsew signal output
rlabel metal2 s 15198 0 15254 800 6 s0_wbd_adr_o[8]
port 349 nsew signal output
rlabel metal2 s 16670 0 16726 800 6 s0_wbd_adr_o[9]
port 350 nsew signal output
rlabel metal2 s 152462 0 152518 800 6 s0_wbd_cyc_o
port 351 nsew signal output
rlabel metal2 s 102874 0 102930 800 6 s0_wbd_dat_i[0]
port 352 nsew signal input
rlabel metal2 s 117410 0 117466 800 6 s0_wbd_dat_i[10]
port 353 nsew signal input
rlabel metal2 s 118882 0 118938 800 6 s0_wbd_dat_i[11]
port 354 nsew signal input
rlabel metal2 s 120354 0 120410 800 6 s0_wbd_dat_i[12]
port 355 nsew signal input
rlabel metal2 s 121826 0 121882 800 6 s0_wbd_dat_i[13]
port 356 nsew signal input
rlabel metal2 s 123298 0 123354 800 6 s0_wbd_dat_i[14]
port 357 nsew signal input
rlabel metal2 s 124770 0 124826 800 6 s0_wbd_dat_i[15]
port 358 nsew signal input
rlabel metal2 s 126242 0 126298 800 6 s0_wbd_dat_i[16]
port 359 nsew signal input
rlabel metal2 s 127622 0 127678 800 6 s0_wbd_dat_i[17]
port 360 nsew signal input
rlabel metal2 s 129094 0 129150 800 6 s0_wbd_dat_i[18]
port 361 nsew signal input
rlabel metal2 s 130566 0 130622 800 6 s0_wbd_dat_i[19]
port 362 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 s0_wbd_dat_i[1]
port 363 nsew signal input
rlabel metal2 s 132038 0 132094 800 6 s0_wbd_dat_i[20]
port 364 nsew signal input
rlabel metal2 s 133510 0 133566 800 6 s0_wbd_dat_i[21]
port 365 nsew signal input
rlabel metal2 s 134982 0 135038 800 6 s0_wbd_dat_i[22]
port 366 nsew signal input
rlabel metal2 s 136454 0 136510 800 6 s0_wbd_dat_i[23]
port 367 nsew signal input
rlabel metal2 s 137926 0 137982 800 6 s0_wbd_dat_i[24]
port 368 nsew signal input
rlabel metal2 s 139306 0 139362 800 6 s0_wbd_dat_i[25]
port 369 nsew signal input
rlabel metal2 s 140778 0 140834 800 6 s0_wbd_dat_i[26]
port 370 nsew signal input
rlabel metal2 s 142250 0 142306 800 6 s0_wbd_dat_i[27]
port 371 nsew signal input
rlabel metal2 s 143722 0 143778 800 6 s0_wbd_dat_i[28]
port 372 nsew signal input
rlabel metal2 s 145194 0 145250 800 6 s0_wbd_dat_i[29]
port 373 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 s0_wbd_dat_i[2]
port 374 nsew signal input
rlabel metal2 s 146666 0 146722 800 6 s0_wbd_dat_i[30]
port 375 nsew signal input
rlabel metal2 s 148138 0 148194 800 6 s0_wbd_dat_i[31]
port 376 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 s0_wbd_dat_i[3]
port 377 nsew signal input
rlabel metal2 s 108670 0 108726 800 6 s0_wbd_dat_i[4]
port 378 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 s0_wbd_dat_i[5]
port 379 nsew signal input
rlabel metal2 s 111614 0 111670 800 6 s0_wbd_dat_i[6]
port 380 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 s0_wbd_dat_i[7]
port 381 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 s0_wbd_dat_i[8]
port 382 nsew signal input
rlabel metal2 s 115938 0 115994 800 6 s0_wbd_dat_i[9]
port 383 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 s0_wbd_dat_o[0]
port 384 nsew signal output
rlabel metal2 s 70674 0 70730 800 6 s0_wbd_dat_o[10]
port 385 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 s0_wbd_dat_o[11]
port 386 nsew signal output
rlabel metal2 s 73618 0 73674 800 6 s0_wbd_dat_o[12]
port 387 nsew signal output
rlabel metal2 s 75090 0 75146 800 6 s0_wbd_dat_o[13]
port 388 nsew signal output
rlabel metal2 s 76562 0 76618 800 6 s0_wbd_dat_o[14]
port 389 nsew signal output
rlabel metal2 s 78034 0 78090 800 6 s0_wbd_dat_o[15]
port 390 nsew signal output
rlabel metal2 s 79506 0 79562 800 6 s0_wbd_dat_o[16]
port 391 nsew signal output
rlabel metal2 s 80978 0 81034 800 6 s0_wbd_dat_o[17]
port 392 nsew signal output
rlabel metal2 s 82358 0 82414 800 6 s0_wbd_dat_o[18]
port 393 nsew signal output
rlabel metal2 s 83830 0 83886 800 6 s0_wbd_dat_o[19]
port 394 nsew signal output
rlabel metal2 s 57610 0 57666 800 6 s0_wbd_dat_o[1]
port 395 nsew signal output
rlabel metal2 s 85302 0 85358 800 6 s0_wbd_dat_o[20]
port 396 nsew signal output
rlabel metal2 s 86774 0 86830 800 6 s0_wbd_dat_o[21]
port 397 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 s0_wbd_dat_o[22]
port 398 nsew signal output
rlabel metal2 s 89718 0 89774 800 6 s0_wbd_dat_o[23]
port 399 nsew signal output
rlabel metal2 s 91190 0 91246 800 6 s0_wbd_dat_o[24]
port 400 nsew signal output
rlabel metal2 s 92662 0 92718 800 6 s0_wbd_dat_o[25]
port 401 nsew signal output
rlabel metal2 s 94042 0 94098 800 6 s0_wbd_dat_o[26]
port 402 nsew signal output
rlabel metal2 s 95514 0 95570 800 6 s0_wbd_dat_o[27]
port 403 nsew signal output
rlabel metal2 s 96986 0 97042 800 6 s0_wbd_dat_o[28]
port 404 nsew signal output
rlabel metal2 s 98458 0 98514 800 6 s0_wbd_dat_o[29]
port 405 nsew signal output
rlabel metal2 s 58990 0 59046 800 6 s0_wbd_dat_o[2]
port 406 nsew signal output
rlabel metal2 s 99930 0 99986 800 6 s0_wbd_dat_o[30]
port 407 nsew signal output
rlabel metal2 s 101402 0 101458 800 6 s0_wbd_dat_o[31]
port 408 nsew signal output
rlabel metal2 s 60462 0 60518 800 6 s0_wbd_dat_o[3]
port 409 nsew signal output
rlabel metal2 s 61934 0 61990 800 6 s0_wbd_dat_o[4]
port 410 nsew signal output
rlabel metal2 s 63406 0 63462 800 6 s0_wbd_dat_o[5]
port 411 nsew signal output
rlabel metal2 s 64878 0 64934 800 6 s0_wbd_dat_o[6]
port 412 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 s0_wbd_dat_o[7]
port 413 nsew signal output
rlabel metal2 s 67822 0 67878 800 6 s0_wbd_dat_o[8]
port 414 nsew signal output
rlabel metal2 s 69294 0 69350 800 6 s0_wbd_dat_o[9]
port 415 nsew signal output
rlabel metal2 s 150990 0 151046 800 6 s0_wbd_err_i
port 416 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 s0_wbd_sel_o[0]
port 417 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 s0_wbd_sel_o[1]
port 418 nsew signal output
rlabel metal2 s 53194 0 53250 800 6 s0_wbd_sel_o[2]
port 419 nsew signal output
rlabel metal2 s 54666 0 54722 800 6 s0_wbd_sel_o[3]
port 420 nsew signal output
rlabel metal2 s 662 0 718 800 6 s0_wbd_stb_o
port 421 nsew signal output
rlabel metal2 s 2042 0 2098 800 6 s0_wbd_we_o
port 422 nsew signal output
rlabel metal2 s 302882 0 302938 800 6 s1_wbd_ack_i
port 423 nsew signal input
rlabel metal2 s 156878 0 156934 800 6 s1_wbd_adr_o[0]
port 424 nsew signal output
rlabel metal2 s 171506 0 171562 800 6 s1_wbd_adr_o[10]
port 425 nsew signal output
rlabel metal2 s 172978 0 173034 800 6 s1_wbd_adr_o[11]
port 426 nsew signal output
rlabel metal2 s 174358 0 174414 800 6 s1_wbd_adr_o[12]
port 427 nsew signal output
rlabel metal2 s 175830 0 175886 800 6 s1_wbd_adr_o[13]
port 428 nsew signal output
rlabel metal2 s 177302 0 177358 800 6 s1_wbd_adr_o[14]
port 429 nsew signal output
rlabel metal2 s 178774 0 178830 800 6 s1_wbd_adr_o[15]
port 430 nsew signal output
rlabel metal2 s 180246 0 180302 800 6 s1_wbd_adr_o[16]
port 431 nsew signal output
rlabel metal2 s 181718 0 181774 800 6 s1_wbd_adr_o[17]
port 432 nsew signal output
rlabel metal2 s 183190 0 183246 800 6 s1_wbd_adr_o[18]
port 433 nsew signal output
rlabel metal2 s 184662 0 184718 800 6 s1_wbd_adr_o[19]
port 434 nsew signal output
rlabel metal2 s 158350 0 158406 800 6 s1_wbd_adr_o[1]
port 435 nsew signal output
rlabel metal2 s 186042 0 186098 800 6 s1_wbd_adr_o[20]
port 436 nsew signal output
rlabel metal2 s 187514 0 187570 800 6 s1_wbd_adr_o[21]
port 437 nsew signal output
rlabel metal2 s 188986 0 189042 800 6 s1_wbd_adr_o[22]
port 438 nsew signal output
rlabel metal2 s 190458 0 190514 800 6 s1_wbd_adr_o[23]
port 439 nsew signal output
rlabel metal2 s 191930 0 191986 800 6 s1_wbd_adr_o[24]
port 440 nsew signal output
rlabel metal2 s 193402 0 193458 800 6 s1_wbd_adr_o[25]
port 441 nsew signal output
rlabel metal2 s 194874 0 194930 800 6 s1_wbd_adr_o[26]
port 442 nsew signal output
rlabel metal2 s 196254 0 196310 800 6 s1_wbd_adr_o[27]
port 443 nsew signal output
rlabel metal2 s 197726 0 197782 800 6 s1_wbd_adr_o[28]
port 444 nsew signal output
rlabel metal2 s 199198 0 199254 800 6 s1_wbd_adr_o[29]
port 445 nsew signal output
rlabel metal2 s 159822 0 159878 800 6 s1_wbd_adr_o[2]
port 446 nsew signal output
rlabel metal2 s 200670 0 200726 800 6 s1_wbd_adr_o[30]
port 447 nsew signal output
rlabel metal2 s 202142 0 202198 800 6 s1_wbd_adr_o[31]
port 448 nsew signal output
rlabel metal2 s 161294 0 161350 800 6 s1_wbd_adr_o[3]
port 449 nsew signal output
rlabel metal2 s 162674 0 162730 800 6 s1_wbd_adr_o[4]
port 450 nsew signal output
rlabel metal2 s 164146 0 164202 800 6 s1_wbd_adr_o[5]
port 451 nsew signal output
rlabel metal2 s 165618 0 165674 800 6 s1_wbd_adr_o[6]
port 452 nsew signal output
rlabel metal2 s 167090 0 167146 800 6 s1_wbd_adr_o[7]
port 453 nsew signal output
rlabel metal2 s 168562 0 168618 800 6 s1_wbd_adr_o[8]
port 454 nsew signal output
rlabel metal2 s 170034 0 170090 800 6 s1_wbd_adr_o[9]
port 455 nsew signal output
rlabel metal2 s 305826 0 305882 800 6 s1_wbd_cyc_o
port 456 nsew signal output
rlabel metal2 s 256146 0 256202 800 6 s1_wbd_dat_i[0]
port 457 nsew signal input
rlabel metal2 s 270774 0 270830 800 6 s1_wbd_dat_i[10]
port 458 nsew signal input
rlabel metal2 s 272246 0 272302 800 6 s1_wbd_dat_i[11]
port 459 nsew signal input
rlabel metal2 s 273718 0 273774 800 6 s1_wbd_dat_i[12]
port 460 nsew signal input
rlabel metal2 s 275190 0 275246 800 6 s1_wbd_dat_i[13]
port 461 nsew signal input
rlabel metal2 s 276662 0 276718 800 6 s1_wbd_dat_i[14]
port 462 nsew signal input
rlabel metal2 s 278042 0 278098 800 6 s1_wbd_dat_i[15]
port 463 nsew signal input
rlabel metal2 s 279514 0 279570 800 6 s1_wbd_dat_i[16]
port 464 nsew signal input
rlabel metal2 s 280986 0 281042 800 6 s1_wbd_dat_i[17]
port 465 nsew signal input
rlabel metal2 s 282458 0 282514 800 6 s1_wbd_dat_i[18]
port 466 nsew signal input
rlabel metal2 s 283930 0 283986 800 6 s1_wbd_dat_i[19]
port 467 nsew signal input
rlabel metal2 s 257618 0 257674 800 6 s1_wbd_dat_i[1]
port 468 nsew signal input
rlabel metal2 s 285402 0 285458 800 6 s1_wbd_dat_i[20]
port 469 nsew signal input
rlabel metal2 s 286874 0 286930 800 6 s1_wbd_dat_i[21]
port 470 nsew signal input
rlabel metal2 s 288254 0 288310 800 6 s1_wbd_dat_i[22]
port 471 nsew signal input
rlabel metal2 s 289726 0 289782 800 6 s1_wbd_dat_i[23]
port 472 nsew signal input
rlabel metal2 s 291198 0 291254 800 6 s1_wbd_dat_i[24]
port 473 nsew signal input
rlabel metal2 s 292670 0 292726 800 6 s1_wbd_dat_i[25]
port 474 nsew signal input
rlabel metal2 s 294142 0 294198 800 6 s1_wbd_dat_i[26]
port 475 nsew signal input
rlabel metal2 s 295614 0 295670 800 6 s1_wbd_dat_i[27]
port 476 nsew signal input
rlabel metal2 s 297086 0 297142 800 6 s1_wbd_dat_i[28]
port 477 nsew signal input
rlabel metal2 s 298558 0 298614 800 6 s1_wbd_dat_i[29]
port 478 nsew signal input
rlabel metal2 s 259090 0 259146 800 6 s1_wbd_dat_i[2]
port 479 nsew signal input
rlabel metal2 s 299938 0 299994 800 6 s1_wbd_dat_i[30]
port 480 nsew signal input
rlabel metal2 s 301410 0 301466 800 6 s1_wbd_dat_i[31]
port 481 nsew signal input
rlabel metal2 s 260562 0 260618 800 6 s1_wbd_dat_i[3]
port 482 nsew signal input
rlabel metal2 s 262034 0 262090 800 6 s1_wbd_dat_i[4]
port 483 nsew signal input
rlabel metal2 s 263506 0 263562 800 6 s1_wbd_dat_i[5]
port 484 nsew signal input
rlabel metal2 s 264978 0 265034 800 6 s1_wbd_dat_i[6]
port 485 nsew signal input
rlabel metal2 s 266358 0 266414 800 6 s1_wbd_dat_i[7]
port 486 nsew signal input
rlabel metal2 s 267830 0 267886 800 6 s1_wbd_dat_i[8]
port 487 nsew signal input
rlabel metal2 s 269302 0 269358 800 6 s1_wbd_dat_i[9]
port 488 nsew signal input
rlabel metal2 s 209410 0 209466 800 6 s1_wbd_dat_o[0]
port 489 nsew signal output
rlabel metal2 s 224038 0 224094 800 6 s1_wbd_dat_o[10]
port 490 nsew signal output
rlabel metal2 s 225510 0 225566 800 6 s1_wbd_dat_o[11]
port 491 nsew signal output
rlabel metal2 s 226982 0 227038 800 6 s1_wbd_dat_o[12]
port 492 nsew signal output
rlabel metal2 s 228454 0 228510 800 6 s1_wbd_dat_o[13]
port 493 nsew signal output
rlabel metal2 s 229926 0 229982 800 6 s1_wbd_dat_o[14]
port 494 nsew signal output
rlabel metal2 s 231306 0 231362 800 6 s1_wbd_dat_o[15]
port 495 nsew signal output
rlabel metal2 s 232778 0 232834 800 6 s1_wbd_dat_o[16]
port 496 nsew signal output
rlabel metal2 s 234250 0 234306 800 6 s1_wbd_dat_o[17]
port 497 nsew signal output
rlabel metal2 s 235722 0 235778 800 6 s1_wbd_dat_o[18]
port 498 nsew signal output
rlabel metal2 s 237194 0 237250 800 6 s1_wbd_dat_o[19]
port 499 nsew signal output
rlabel metal2 s 210882 0 210938 800 6 s1_wbd_dat_o[1]
port 500 nsew signal output
rlabel metal2 s 238666 0 238722 800 6 s1_wbd_dat_o[20]
port 501 nsew signal output
rlabel metal2 s 240138 0 240194 800 6 s1_wbd_dat_o[21]
port 502 nsew signal output
rlabel metal2 s 241610 0 241666 800 6 s1_wbd_dat_o[22]
port 503 nsew signal output
rlabel metal2 s 242990 0 243046 800 6 s1_wbd_dat_o[23]
port 504 nsew signal output
rlabel metal2 s 244462 0 244518 800 6 s1_wbd_dat_o[24]
port 505 nsew signal output
rlabel metal2 s 245934 0 245990 800 6 s1_wbd_dat_o[25]
port 506 nsew signal output
rlabel metal2 s 247406 0 247462 800 6 s1_wbd_dat_o[26]
port 507 nsew signal output
rlabel metal2 s 248878 0 248934 800 6 s1_wbd_dat_o[27]
port 508 nsew signal output
rlabel metal2 s 250350 0 250406 800 6 s1_wbd_dat_o[28]
port 509 nsew signal output
rlabel metal2 s 251822 0 251878 800 6 s1_wbd_dat_o[29]
port 510 nsew signal output
rlabel metal2 s 212354 0 212410 800 6 s1_wbd_dat_o[2]
port 511 nsew signal output
rlabel metal2 s 253294 0 253350 800 6 s1_wbd_dat_o[30]
port 512 nsew signal output
rlabel metal2 s 254674 0 254730 800 6 s1_wbd_dat_o[31]
port 513 nsew signal output
rlabel metal2 s 213826 0 213882 800 6 s1_wbd_dat_o[3]
port 514 nsew signal output
rlabel metal2 s 215298 0 215354 800 6 s1_wbd_dat_o[4]
port 515 nsew signal output
rlabel metal2 s 216770 0 216826 800 6 s1_wbd_dat_o[5]
port 516 nsew signal output
rlabel metal2 s 218242 0 218298 800 6 s1_wbd_dat_o[6]
port 517 nsew signal output
rlabel metal2 s 219622 0 219678 800 6 s1_wbd_dat_o[7]
port 518 nsew signal output
rlabel metal2 s 221094 0 221150 800 6 s1_wbd_dat_o[8]
port 519 nsew signal output
rlabel metal2 s 222566 0 222622 800 6 s1_wbd_dat_o[9]
port 520 nsew signal output
rlabel metal2 s 304354 0 304410 800 6 s1_wbd_err_i
port 521 nsew signal input
rlabel metal2 s 203614 0 203670 800 6 s1_wbd_sel_o[0]
port 522 nsew signal output
rlabel metal2 s 205086 0 205142 800 6 s1_wbd_sel_o[1]
port 523 nsew signal output
rlabel metal2 s 206558 0 206614 800 6 s1_wbd_sel_o[2]
port 524 nsew signal output
rlabel metal2 s 207938 0 207994 800 6 s1_wbd_sel_o[3]
port 525 nsew signal output
rlabel metal2 s 153934 0 153990 800 6 s1_wbd_stb_o
port 526 nsew signal output
rlabel metal2 s 155406 0 155462 800 6 s1_wbd_we_o
port 527 nsew signal output
rlabel metal2 s 456246 0 456302 800 6 s2_wbd_ack_i
port 528 nsew signal input
rlabel metal2 s 310242 0 310298 800 6 s2_wbd_adr_o[0]
port 529 nsew signal output
rlabel metal2 s 324778 0 324834 800 6 s2_wbd_adr_o[10]
port 530 nsew signal output
rlabel metal2 s 326250 0 326306 800 6 s2_wbd_adr_o[11]
port 531 nsew signal output
rlabel metal2 s 327722 0 327778 800 6 s2_wbd_adr_o[12]
port 532 nsew signal output
rlabel metal2 s 329194 0 329250 800 6 s2_wbd_adr_o[13]
port 533 nsew signal output
rlabel metal2 s 330666 0 330722 800 6 s2_wbd_adr_o[14]
port 534 nsew signal output
rlabel metal2 s 332138 0 332194 800 6 s2_wbd_adr_o[15]
port 535 nsew signal output
rlabel metal2 s 333610 0 333666 800 6 s2_wbd_adr_o[16]
port 536 nsew signal output
rlabel metal2 s 334990 0 335046 800 6 s2_wbd_adr_o[17]
port 537 nsew signal output
rlabel metal2 s 336462 0 336518 800 6 s2_wbd_adr_o[18]
port 538 nsew signal output
rlabel metal2 s 337934 0 337990 800 6 s2_wbd_adr_o[19]
port 539 nsew signal output
rlabel metal2 s 311622 0 311678 800 6 s2_wbd_adr_o[1]
port 540 nsew signal output
rlabel metal2 s 339406 0 339462 800 6 s2_wbd_adr_o[20]
port 541 nsew signal output
rlabel metal2 s 340878 0 340934 800 6 s2_wbd_adr_o[21]
port 542 nsew signal output
rlabel metal2 s 342350 0 342406 800 6 s2_wbd_adr_o[22]
port 543 nsew signal output
rlabel metal2 s 343822 0 343878 800 6 s2_wbd_adr_o[23]
port 544 nsew signal output
rlabel metal2 s 345294 0 345350 800 6 s2_wbd_adr_o[24]
port 545 nsew signal output
rlabel metal2 s 346674 0 346730 800 6 s2_wbd_adr_o[25]
port 546 nsew signal output
rlabel metal2 s 348146 0 348202 800 6 s2_wbd_adr_o[26]
port 547 nsew signal output
rlabel metal2 s 349618 0 349674 800 6 s2_wbd_adr_o[27]
port 548 nsew signal output
rlabel metal2 s 351090 0 351146 800 6 s2_wbd_adr_o[28]
port 549 nsew signal output
rlabel metal2 s 352562 0 352618 800 6 s2_wbd_adr_o[29]
port 550 nsew signal output
rlabel metal2 s 313094 0 313150 800 6 s2_wbd_adr_o[2]
port 551 nsew signal output
rlabel metal2 s 354034 0 354090 800 6 s2_wbd_adr_o[30]
port 552 nsew signal output
rlabel metal2 s 355506 0 355562 800 6 s2_wbd_adr_o[31]
port 553 nsew signal output
rlabel metal2 s 314566 0 314622 800 6 s2_wbd_adr_o[3]
port 554 nsew signal output
rlabel metal2 s 316038 0 316094 800 6 s2_wbd_adr_o[4]
port 555 nsew signal output
rlabel metal2 s 317510 0 317566 800 6 s2_wbd_adr_o[5]
port 556 nsew signal output
rlabel metal2 s 318982 0 319038 800 6 s2_wbd_adr_o[6]
port 557 nsew signal output
rlabel metal2 s 320454 0 320510 800 6 s2_wbd_adr_o[7]
port 558 nsew signal output
rlabel metal2 s 321926 0 321982 800 6 s2_wbd_adr_o[8]
port 559 nsew signal output
rlabel metal2 s 323306 0 323362 800 6 s2_wbd_adr_o[9]
port 560 nsew signal output
rlabel metal2 s 459190 0 459246 800 6 s2_wbd_cyc_o
port 561 nsew signal output
rlabel metal2 s 409510 0 409566 800 6 s2_wbd_dat_i[0]
port 562 nsew signal input
rlabel metal2 s 424138 0 424194 800 6 s2_wbd_dat_i[10]
port 563 nsew signal input
rlabel metal2 s 425610 0 425666 800 6 s2_wbd_dat_i[11]
port 564 nsew signal input
rlabel metal2 s 426990 0 427046 800 6 s2_wbd_dat_i[12]
port 565 nsew signal input
rlabel metal2 s 428462 0 428518 800 6 s2_wbd_dat_i[13]
port 566 nsew signal input
rlabel metal2 s 429934 0 429990 800 6 s2_wbd_dat_i[14]
port 567 nsew signal input
rlabel metal2 s 431406 0 431462 800 6 s2_wbd_dat_i[15]
port 568 nsew signal input
rlabel metal2 s 432878 0 432934 800 6 s2_wbd_dat_i[16]
port 569 nsew signal input
rlabel metal2 s 434350 0 434406 800 6 s2_wbd_dat_i[17]
port 570 nsew signal input
rlabel metal2 s 435822 0 435878 800 6 s2_wbd_dat_i[18]
port 571 nsew signal input
rlabel metal2 s 437294 0 437350 800 6 s2_wbd_dat_i[19]
port 572 nsew signal input
rlabel metal2 s 410982 0 411038 800 6 s2_wbd_dat_i[1]
port 573 nsew signal input
rlabel metal2 s 438674 0 438730 800 6 s2_wbd_dat_i[20]
port 574 nsew signal input
rlabel metal2 s 440146 0 440202 800 6 s2_wbd_dat_i[21]
port 575 nsew signal input
rlabel metal2 s 441618 0 441674 800 6 s2_wbd_dat_i[22]
port 576 nsew signal input
rlabel metal2 s 443090 0 443146 800 6 s2_wbd_dat_i[23]
port 577 nsew signal input
rlabel metal2 s 444562 0 444618 800 6 s2_wbd_dat_i[24]
port 578 nsew signal input
rlabel metal2 s 446034 0 446090 800 6 s2_wbd_dat_i[25]
port 579 nsew signal input
rlabel metal2 s 447506 0 447562 800 6 s2_wbd_dat_i[26]
port 580 nsew signal input
rlabel metal2 s 448978 0 449034 800 6 s2_wbd_dat_i[27]
port 581 nsew signal input
rlabel metal2 s 450358 0 450414 800 6 s2_wbd_dat_i[28]
port 582 nsew signal input
rlabel metal2 s 451830 0 451886 800 6 s2_wbd_dat_i[29]
port 583 nsew signal input
rlabel metal2 s 412454 0 412510 800 6 s2_wbd_dat_i[2]
port 584 nsew signal input
rlabel metal2 s 453302 0 453358 800 6 s2_wbd_dat_i[30]
port 585 nsew signal input
rlabel metal2 s 454774 0 454830 800 6 s2_wbd_dat_i[31]
port 586 nsew signal input
rlabel metal2 s 413926 0 413982 800 6 s2_wbd_dat_i[3]
port 587 nsew signal input
rlabel metal2 s 415306 0 415362 800 6 s2_wbd_dat_i[4]
port 588 nsew signal input
rlabel metal2 s 416778 0 416834 800 6 s2_wbd_dat_i[5]
port 589 nsew signal input
rlabel metal2 s 418250 0 418306 800 6 s2_wbd_dat_i[6]
port 590 nsew signal input
rlabel metal2 s 419722 0 419778 800 6 s2_wbd_dat_i[7]
port 591 nsew signal input
rlabel metal2 s 421194 0 421250 800 6 s2_wbd_dat_i[8]
port 592 nsew signal input
rlabel metal2 s 422666 0 422722 800 6 s2_wbd_dat_i[9]
port 593 nsew signal input
rlabel metal2 s 362774 0 362830 800 6 s2_wbd_dat_o[0]
port 594 nsew signal output
rlabel metal2 s 377402 0 377458 800 6 s2_wbd_dat_o[10]
port 595 nsew signal output
rlabel metal2 s 378874 0 378930 800 6 s2_wbd_dat_o[11]
port 596 nsew signal output
rlabel metal2 s 380254 0 380310 800 6 s2_wbd_dat_o[12]
port 597 nsew signal output
rlabel metal2 s 381726 0 381782 800 6 s2_wbd_dat_o[13]
port 598 nsew signal output
rlabel metal2 s 383198 0 383254 800 6 s2_wbd_dat_o[14]
port 599 nsew signal output
rlabel metal2 s 384670 0 384726 800 6 s2_wbd_dat_o[15]
port 600 nsew signal output
rlabel metal2 s 386142 0 386198 800 6 s2_wbd_dat_o[16]
port 601 nsew signal output
rlabel metal2 s 387614 0 387670 800 6 s2_wbd_dat_o[17]
port 602 nsew signal output
rlabel metal2 s 389086 0 389142 800 6 s2_wbd_dat_o[18]
port 603 nsew signal output
rlabel metal2 s 390558 0 390614 800 6 s2_wbd_dat_o[19]
port 604 nsew signal output
rlabel metal2 s 364246 0 364302 800 6 s2_wbd_dat_o[1]
port 605 nsew signal output
rlabel metal2 s 391938 0 391994 800 6 s2_wbd_dat_o[20]
port 606 nsew signal output
rlabel metal2 s 393410 0 393466 800 6 s2_wbd_dat_o[21]
port 607 nsew signal output
rlabel metal2 s 394882 0 394938 800 6 s2_wbd_dat_o[22]
port 608 nsew signal output
rlabel metal2 s 396354 0 396410 800 6 s2_wbd_dat_o[23]
port 609 nsew signal output
rlabel metal2 s 397826 0 397882 800 6 s2_wbd_dat_o[24]
port 610 nsew signal output
rlabel metal2 s 399298 0 399354 800 6 s2_wbd_dat_o[25]
port 611 nsew signal output
rlabel metal2 s 400770 0 400826 800 6 s2_wbd_dat_o[26]
port 612 nsew signal output
rlabel metal2 s 402242 0 402298 800 6 s2_wbd_dat_o[27]
port 613 nsew signal output
rlabel metal2 s 403622 0 403678 800 6 s2_wbd_dat_o[28]
port 614 nsew signal output
rlabel metal2 s 405094 0 405150 800 6 s2_wbd_dat_o[29]
port 615 nsew signal output
rlabel metal2 s 365718 0 365774 800 6 s2_wbd_dat_o[2]
port 616 nsew signal output
rlabel metal2 s 406566 0 406622 800 6 s2_wbd_dat_o[30]
port 617 nsew signal output
rlabel metal2 s 408038 0 408094 800 6 s2_wbd_dat_o[31]
port 618 nsew signal output
rlabel metal2 s 367190 0 367246 800 6 s2_wbd_dat_o[3]
port 619 nsew signal output
rlabel metal2 s 368662 0 368718 800 6 s2_wbd_dat_o[4]
port 620 nsew signal output
rlabel metal2 s 370042 0 370098 800 6 s2_wbd_dat_o[5]
port 621 nsew signal output
rlabel metal2 s 371514 0 371570 800 6 s2_wbd_dat_o[6]
port 622 nsew signal output
rlabel metal2 s 372986 0 373042 800 6 s2_wbd_dat_o[7]
port 623 nsew signal output
rlabel metal2 s 374458 0 374514 800 6 s2_wbd_dat_o[8]
port 624 nsew signal output
rlabel metal2 s 375930 0 375986 800 6 s2_wbd_dat_o[9]
port 625 nsew signal output
rlabel metal2 s 457718 0 457774 800 6 s2_wbd_err_i
port 626 nsew signal input
rlabel metal2 s 356978 0 357034 800 6 s2_wbd_sel_o[0]
port 627 nsew signal output
rlabel metal2 s 358358 0 358414 800 6 s2_wbd_sel_o[1]
port 628 nsew signal output
rlabel metal2 s 359830 0 359886 800 6 s2_wbd_sel_o[2]
port 629 nsew signal output
rlabel metal2 s 361302 0 361358 800 6 s2_wbd_sel_o[3]
port 630 nsew signal output
rlabel metal2 s 307298 0 307354 800 6 s2_wbd_stb_o
port 631 nsew signal output
rlabel metal2 s 308770 0 308826 800 6 s2_wbd_we_o
port 632 nsew signal output
rlabel metal2 s 451350 1040 451410 18544 6 VPWR
port 633 nsew power bidirectional
rlabel metal2 s 435350 1040 435410 18544 6 VPWR
port 634 nsew power bidirectional
rlabel metal2 s 419350 1040 419410 18544 6 VPWR
port 635 nsew power bidirectional
rlabel metal2 s 403350 1040 403410 18544 6 VPWR
port 636 nsew power bidirectional
rlabel metal2 s 387350 1040 387410 18544 6 VPWR
port 637 nsew power bidirectional
rlabel metal2 s 371350 1040 371410 18544 6 VPWR
port 638 nsew power bidirectional
rlabel metal2 s 355350 1040 355410 18544 6 VPWR
port 639 nsew power bidirectional
rlabel metal2 s 339350 1040 339410 18544 6 VPWR
port 640 nsew power bidirectional
rlabel metal2 s 323350 1040 323410 18544 6 VPWR
port 641 nsew power bidirectional
rlabel metal2 s 307350 1040 307410 18544 6 VPWR
port 642 nsew power bidirectional
rlabel metal2 s 291350 1040 291410 18544 6 VPWR
port 643 nsew power bidirectional
rlabel metal2 s 275350 1040 275410 18544 6 VPWR
port 644 nsew power bidirectional
rlabel metal2 s 259350 1040 259410 18544 6 VPWR
port 645 nsew power bidirectional
rlabel metal2 s 243350 1040 243410 18544 6 VPWR
port 646 nsew power bidirectional
rlabel metal2 s 227350 1040 227410 18544 6 VPWR
port 647 nsew power bidirectional
rlabel metal2 s 211350 1040 211410 18544 6 VPWR
port 648 nsew power bidirectional
rlabel metal2 s 195350 1040 195410 18544 6 VPWR
port 649 nsew power bidirectional
rlabel metal2 s 179350 1040 179410 18544 6 VPWR
port 650 nsew power bidirectional
rlabel metal2 s 163350 1040 163410 18544 6 VPWR
port 651 nsew power bidirectional
rlabel metal2 s 147350 1040 147410 18544 6 VPWR
port 652 nsew power bidirectional
rlabel metal2 s 131350 1040 131410 18544 6 VPWR
port 653 nsew power bidirectional
rlabel metal2 s 115350 1040 115410 18544 6 VPWR
port 654 nsew power bidirectional
rlabel metal2 s 99350 1040 99410 18544 6 VPWR
port 655 nsew power bidirectional
rlabel metal2 s 83350 1040 83410 18544 6 VPWR
port 656 nsew power bidirectional
rlabel metal2 s 67350 1040 67410 18544 6 VPWR
port 657 nsew power bidirectional
rlabel metal2 s 51350 1040 51410 18544 6 VPWR
port 658 nsew power bidirectional
rlabel metal2 s 35350 1040 35410 18544 6 VPWR
port 659 nsew power bidirectional
rlabel metal2 s 19350 1040 19410 18544 6 VPWR
port 660 nsew power bidirectional
rlabel metal2 s 3350 1040 3410 18544 6 VPWR
port 661 nsew power bidirectional
rlabel metal3 s 1380 16330 458620 16390 6 VPWR
port 662 nsew power bidirectional
rlabel metal3 s 1380 14170 458620 14230 6 VPWR
port 663 nsew power bidirectional
rlabel metal3 s 1380 12010 458620 12070 6 VPWR
port 664 nsew power bidirectional
rlabel metal3 s 1380 9850 458620 9910 6 VPWR
port 665 nsew power bidirectional
rlabel metal3 s 1380 7690 458620 7750 6 VPWR
port 666 nsew power bidirectional
rlabel metal3 s 1380 5530 458620 5590 6 VPWR
port 667 nsew power bidirectional
rlabel metal3 s 1380 3370 458620 3430 6 VPWR
port 668 nsew power bidirectional
rlabel metal3 s 1380 1210 458620 1270 6 VPWR
port 669 nsew power bidirectional
rlabel metal2 s 443350 1040 443410 18544 6 VGND
port 670 nsew ground bidirectional
rlabel metal2 s 427350 1040 427410 18544 6 VGND
port 671 nsew ground bidirectional
rlabel metal2 s 411350 1040 411410 18544 6 VGND
port 672 nsew ground bidirectional
rlabel metal2 s 395350 1040 395410 18544 6 VGND
port 673 nsew ground bidirectional
rlabel metal2 s 379350 1040 379410 18544 6 VGND
port 674 nsew ground bidirectional
rlabel metal2 s 363350 1040 363410 18544 6 VGND
port 675 nsew ground bidirectional
rlabel metal2 s 347350 1040 347410 18544 6 VGND
port 676 nsew ground bidirectional
rlabel metal2 s 331350 1040 331410 18544 6 VGND
port 677 nsew ground bidirectional
rlabel metal2 s 315350 1040 315410 18544 6 VGND
port 678 nsew ground bidirectional
rlabel metal2 s 299350 1040 299410 18544 6 VGND
port 679 nsew ground bidirectional
rlabel metal2 s 283350 1040 283410 18544 6 VGND
port 680 nsew ground bidirectional
rlabel metal2 s 267350 1040 267410 18544 6 VGND
port 681 nsew ground bidirectional
rlabel metal2 s 251350 1040 251410 18544 6 VGND
port 682 nsew ground bidirectional
rlabel metal2 s 235350 1040 235410 18544 6 VGND
port 683 nsew ground bidirectional
rlabel metal2 s 219350 1040 219410 18544 6 VGND
port 684 nsew ground bidirectional
rlabel metal2 s 203350 1040 203410 18544 6 VGND
port 685 nsew ground bidirectional
rlabel metal2 s 187350 1040 187410 18544 6 VGND
port 686 nsew ground bidirectional
rlabel metal2 s 171350 1040 171410 18544 6 VGND
port 687 nsew ground bidirectional
rlabel metal2 s 155350 1040 155410 18544 6 VGND
port 688 nsew ground bidirectional
rlabel metal2 s 139350 1040 139410 18544 6 VGND
port 689 nsew ground bidirectional
rlabel metal2 s 123350 1040 123410 18544 6 VGND
port 690 nsew ground bidirectional
rlabel metal2 s 107350 1040 107410 18544 6 VGND
port 691 nsew ground bidirectional
rlabel metal2 s 91350 1040 91410 18544 6 VGND
port 692 nsew ground bidirectional
rlabel metal2 s 75350 1040 75410 18544 6 VGND
port 693 nsew ground bidirectional
rlabel metal2 s 59350 1040 59410 18544 6 VGND
port 694 nsew ground bidirectional
rlabel metal2 s 43350 1040 43410 18544 6 VGND
port 695 nsew ground bidirectional
rlabel metal2 s 27350 1040 27410 18544 6 VGND
port 696 nsew ground bidirectional
rlabel metal2 s 11350 1040 11410 18544 6 VGND
port 697 nsew ground bidirectional
rlabel metal3 s 1380 17410 458620 17470 6 VGND
port 698 nsew ground bidirectional
rlabel metal3 s 1380 15250 458620 15310 6 VGND
port 699 nsew ground bidirectional
rlabel metal3 s 1380 13090 458620 13150 6 VGND
port 700 nsew ground bidirectional
rlabel metal3 s 1380 10930 458620 10990 6 VGND
port 701 nsew ground bidirectional
rlabel metal3 s 1380 8770 458620 8830 6 VGND
port 702 nsew ground bidirectional
rlabel metal3 s 1380 6610 458620 6670 6 VGND
port 703 nsew ground bidirectional
rlabel metal3 s 1380 4450 458620 4510 6 VGND
port 704 nsew ground bidirectional
rlabel metal3 s 1380 2290 458620 2350 6 VGND
port 705 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 460000 20000
string LEFview TRUE
string GDS_FILE /project/openlane/wb_interconnect/runs/wb_interconnect/results/magic/wb_interconnect.gds
string GDS_END 5210272
string GDS_START 199828
<< end >>

