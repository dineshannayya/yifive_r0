magic
tech sky130A
magscale 1 2
timestamp 1623923575
<< obsli1 >>
rect 1380 1071 58604 58769
<< obsm1 >>
rect 382 892 59602 59016
<< metal2 >>
rect 386 59200 442 60000
rect 1122 59200 1178 60000
rect 1950 59200 2006 60000
rect 2686 59200 2742 60000
rect 3514 59200 3570 60000
rect 4250 59200 4306 60000
rect 5078 59200 5134 60000
rect 5906 59200 5962 60000
rect 6642 59200 6698 60000
rect 7470 59200 7526 60000
rect 8206 59200 8262 60000
rect 9034 59200 9090 60000
rect 9770 59200 9826 60000
rect 10598 59200 10654 60000
rect 11426 59200 11482 60000
rect 12162 59200 12218 60000
rect 12990 59200 13046 60000
rect 13726 59200 13782 60000
rect 14554 59200 14610 60000
rect 15382 59200 15438 60000
rect 16118 59200 16174 60000
rect 16946 59200 17002 60000
rect 17682 59200 17738 60000
rect 18510 59200 18566 60000
rect 19246 59200 19302 60000
rect 20074 59200 20130 60000
rect 20902 59200 20958 60000
rect 21638 59200 21694 60000
rect 22466 59200 22522 60000
rect 23202 59200 23258 60000
rect 24030 59200 24086 60000
rect 24766 59200 24822 60000
rect 25594 59200 25650 60000
rect 26422 59200 26478 60000
rect 27158 59200 27214 60000
rect 27986 59200 28042 60000
rect 28722 59200 28778 60000
rect 29550 59200 29606 60000
rect 30378 59200 30434 60000
rect 31114 59200 31170 60000
rect 31942 59200 31998 60000
rect 32678 59200 32734 60000
rect 33506 59200 33562 60000
rect 34242 59200 34298 60000
rect 35070 59200 35126 60000
rect 35898 59200 35954 60000
rect 36634 59200 36690 60000
rect 37462 59200 37518 60000
rect 38198 59200 38254 60000
rect 39026 59200 39082 60000
rect 39762 59200 39818 60000
rect 40590 59200 40646 60000
rect 41418 59200 41474 60000
rect 42154 59200 42210 60000
rect 42982 59200 43038 60000
rect 43718 59200 43774 60000
rect 44546 59200 44602 60000
rect 45374 59200 45430 60000
rect 46110 59200 46166 60000
rect 46938 59200 46994 60000
rect 47674 59200 47730 60000
rect 48502 59200 48558 60000
rect 49238 59200 49294 60000
rect 50066 59200 50122 60000
rect 50894 59200 50950 60000
rect 51630 59200 51686 60000
rect 52458 59200 52514 60000
rect 53194 59200 53250 60000
rect 54022 59200 54078 60000
rect 54758 59200 54814 60000
rect 55586 59200 55642 60000
rect 56414 59200 56470 60000
rect 57150 59200 57206 60000
rect 57978 59200 58034 60000
rect 58714 59200 58770 60000
rect 59542 59200 59598 60000
rect 3350 1040 3410 58800
rect 11350 1040 11410 58800
rect 19350 1040 19410 58800
rect 27350 1040 27410 58800
rect 35350 1040 35410 58800
rect 43350 1040 43410 58800
rect 51350 1040 51410 58800
rect 30010 0 30066 800
<< obsm2 >>
rect 498 59144 1066 59537
rect 1234 59144 1894 59537
rect 2062 59144 2630 59537
rect 2798 59144 3458 59537
rect 3626 59144 4194 59537
rect 4362 59144 5022 59537
rect 5190 59144 5850 59537
rect 6018 59144 6586 59537
rect 6754 59144 7414 59537
rect 7582 59144 8150 59537
rect 8318 59144 8978 59537
rect 9146 59144 9714 59537
rect 9882 59144 10542 59537
rect 10710 59144 11370 59537
rect 11538 59144 12106 59537
rect 12274 59144 12934 59537
rect 13102 59144 13670 59537
rect 13838 59144 14498 59537
rect 14666 59144 15326 59537
rect 15494 59144 16062 59537
rect 16230 59144 16890 59537
rect 17058 59144 17626 59537
rect 17794 59144 18454 59537
rect 18622 59144 19190 59537
rect 19358 59144 20018 59537
rect 20186 59144 20846 59537
rect 21014 59144 21582 59537
rect 21750 59144 22410 59537
rect 22578 59144 23146 59537
rect 23314 59144 23974 59537
rect 24142 59144 24710 59537
rect 24878 59144 25538 59537
rect 25706 59144 26366 59537
rect 26534 59144 27102 59537
rect 27270 59144 27930 59537
rect 28098 59144 28666 59537
rect 28834 59144 29494 59537
rect 29662 59144 30322 59537
rect 30490 59144 31058 59537
rect 31226 59144 31886 59537
rect 32054 59144 32622 59537
rect 32790 59144 33450 59537
rect 33618 59144 34186 59537
rect 34354 59144 35014 59537
rect 35182 59144 35842 59537
rect 36010 59144 36578 59537
rect 36746 59144 37406 59537
rect 37574 59144 38142 59537
rect 38310 59144 38970 59537
rect 39138 59144 39706 59537
rect 39874 59144 40534 59537
rect 40702 59144 41362 59537
rect 41530 59144 42098 59537
rect 42266 59144 42926 59537
rect 43094 59144 43662 59537
rect 43830 59144 44490 59537
rect 44658 59144 45318 59537
rect 45486 59144 46054 59537
rect 46222 59144 46882 59537
rect 47050 59144 47618 59537
rect 47786 59144 48446 59537
rect 48614 59144 49182 59537
rect 49350 59144 50010 59537
rect 50178 59144 50838 59537
rect 51006 59144 51574 59537
rect 51742 59144 52402 59537
rect 52570 59144 53138 59537
rect 53306 59144 53966 59537
rect 54134 59144 54702 59537
rect 54870 59144 55530 59537
rect 55698 59144 56358 59537
rect 56526 59144 57094 59537
rect 57262 59144 57922 59537
rect 58090 59144 58658 59537
rect 58826 59144 59486 59537
rect 388 58856 59596 59144
rect 388 984 3294 58856
rect 3466 984 11294 58856
rect 11466 984 19294 58856
rect 19466 984 27294 58856
rect 27466 984 35294 58856
rect 35466 984 43294 58856
rect 43466 984 51294 58856
rect 51466 984 59596 58856
rect 388 856 59596 984
rect 388 303 29954 856
rect 30122 303 59596 856
<< metal3 >>
rect 0 59304 800 59424
rect 59200 59440 60000 59560
rect 59200 58760 60000 58880
rect 0 58352 800 58472
rect 1380 58450 58604 58510
rect 59200 58080 60000 58200
rect 0 57400 800 57520
rect 1380 57370 58604 57430
rect 59200 57400 60000 57520
rect 59200 56720 60000 56840
rect 0 56448 800 56568
rect 1380 56290 58604 56350
rect 59200 56040 60000 56160
rect 0 55360 800 55480
rect 59200 55360 60000 55480
rect 1380 55210 58604 55270
rect 0 54408 800 54528
rect 59200 54544 60000 54664
rect 1380 54130 58604 54190
rect 59200 53864 60000 53984
rect 0 53456 800 53576
rect 1380 53050 58604 53110
rect 59200 53184 60000 53304
rect 0 52504 800 52624
rect 59200 52504 60000 52624
rect 1380 51970 58604 52030
rect 59200 51824 60000 51944
rect 0 51416 800 51536
rect 59200 51144 60000 51264
rect 1380 50890 58604 50950
rect 0 50464 800 50584
rect 59200 50464 60000 50584
rect 1380 49810 58604 49870
rect 59200 49784 60000 49904
rect 0 49512 800 49632
rect 59200 48968 60000 49088
rect 0 48560 800 48680
rect 1380 48730 58604 48790
rect 59200 48288 60000 48408
rect 0 47608 800 47728
rect 1380 47650 58604 47710
rect 59200 47608 60000 47728
rect 59200 46928 60000 47048
rect 0 46520 800 46640
rect 1380 46570 58604 46630
rect 59200 46248 60000 46368
rect 0 45568 800 45688
rect 1380 45490 58604 45550
rect 59200 45568 60000 45688
rect 59200 44888 60000 45008
rect 0 44616 800 44736
rect 1380 44410 58604 44470
rect 59200 44208 60000 44328
rect 0 43664 800 43784
rect 1380 43330 58604 43390
rect 59200 43392 60000 43512
rect 0 42576 800 42696
rect 59200 42712 60000 42832
rect 1380 42250 58604 42310
rect 59200 42032 60000 42152
rect 0 41624 800 41744
rect 59200 41352 60000 41472
rect 1380 41170 58604 41230
rect 0 40672 800 40792
rect 59200 40672 60000 40792
rect 1380 40090 58604 40150
rect 59200 39992 60000 40112
rect 0 39720 800 39840
rect 59200 39312 60000 39432
rect 1380 39010 58604 39070
rect 0 38632 800 38752
rect 59200 38632 60000 38752
rect 1380 37930 58604 37990
rect 0 37680 800 37800
rect 59200 37816 60000 37936
rect 59200 37136 60000 37256
rect 0 36728 800 36848
rect 1380 36850 58604 36910
rect 59200 36456 60000 36576
rect 0 35776 800 35896
rect 1380 35770 58604 35830
rect 59200 35776 60000 35896
rect 59200 35096 60000 35216
rect 0 34824 800 34944
rect 1380 34690 58604 34750
rect 59200 34416 60000 34536
rect 0 33736 800 33856
rect 1380 33610 58604 33670
rect 59200 33736 60000 33856
rect 59200 33056 60000 33176
rect 0 32784 800 32904
rect 1380 32530 58604 32590
rect 59200 32240 60000 32360
rect 0 31832 800 31952
rect 1380 31450 58604 31510
rect 59200 31560 60000 31680
rect 0 30880 800 31000
rect 59200 30880 60000 31000
rect 1380 30370 58604 30430
rect 59200 30200 60000 30320
rect 0 29792 800 29912
rect 59200 29520 60000 29640
rect 1380 29290 58604 29350
rect 0 28840 800 28960
rect 59200 28840 60000 28960
rect 1380 28210 58604 28270
rect 59200 28160 60000 28280
rect 0 27888 800 28008
rect 59200 27344 60000 27464
rect 0 26936 800 27056
rect 1380 27130 58604 27190
rect 59200 26664 60000 26784
rect 1380 26050 58604 26110
rect 59200 25984 60000 26104
rect 0 25848 800 25968
rect 59200 25304 60000 25424
rect 0 24896 800 25016
rect 1380 24970 58604 25030
rect 59200 24624 60000 24744
rect 0 23944 800 24064
rect 1380 23890 58604 23950
rect 59200 23944 60000 24064
rect 59200 23264 60000 23384
rect 0 22992 800 23112
rect 1380 22810 58604 22870
rect 59200 22584 60000 22704
rect 0 22040 800 22160
rect 1380 21730 58604 21790
rect 59200 21768 60000 21888
rect 0 20952 800 21072
rect 59200 21088 60000 21208
rect 1380 20650 58604 20710
rect 59200 20408 60000 20528
rect 0 20000 800 20120
rect 59200 19728 60000 19848
rect 1380 19570 58604 19630
rect 0 19048 800 19168
rect 59200 19048 60000 19168
rect 1380 18490 58604 18550
rect 59200 18368 60000 18488
rect 0 18096 800 18216
rect 59200 17688 60000 17808
rect 1380 17410 58604 17470
rect 0 17008 800 17128
rect 59200 17008 60000 17128
rect 1380 16330 58604 16390
rect 0 16056 800 16176
rect 59200 16192 60000 16312
rect 59200 15512 60000 15632
rect 0 15104 800 15224
rect 1380 15250 58604 15310
rect 59200 14832 60000 14952
rect 0 14152 800 14272
rect 1380 14170 58604 14230
rect 59200 14152 60000 14272
rect 59200 13472 60000 13592
rect 0 13064 800 13184
rect 1380 13090 58604 13150
rect 59200 12792 60000 12912
rect 0 12112 800 12232
rect 1380 12010 58604 12070
rect 59200 12112 60000 12232
rect 59200 11432 60000 11552
rect 0 11160 800 11280
rect 1380 10930 58604 10990
rect 59200 10616 60000 10736
rect 0 10208 800 10328
rect 1380 9850 58604 9910
rect 59200 9936 60000 10056
rect 0 9256 800 9376
rect 59200 9256 60000 9376
rect 1380 8770 58604 8830
rect 59200 8576 60000 8696
rect 0 8168 800 8288
rect 59200 7896 60000 8016
rect 1380 7690 58604 7750
rect 0 7216 800 7336
rect 59200 7216 60000 7336
rect 1380 6610 58604 6670
rect 59200 6536 60000 6656
rect 0 6264 800 6384
rect 59200 5856 60000 5976
rect 1380 5530 58604 5590
rect 0 5312 800 5432
rect 59200 5040 60000 5160
rect 1380 4450 58604 4510
rect 0 4224 800 4344
rect 59200 4360 60000 4480
rect 59200 3680 60000 3800
rect 0 3272 800 3392
rect 1380 3370 58604 3430
rect 59200 3000 60000 3120
rect 0 2320 800 2440
rect 1380 2290 58604 2350
rect 59200 2320 60000 2440
rect 59200 1640 60000 1760
rect 0 1368 800 1488
rect 1380 1210 58604 1270
rect 59200 960 60000 1080
rect 0 416 800 536
rect 59200 280 60000 400
<< obsm3 >>
rect 800 59504 59120 59533
rect 880 59360 59120 59504
rect 880 59224 59200 59360
rect 800 58960 59200 59224
rect 800 58680 59120 58960
rect 800 58590 59200 58680
rect 800 58552 1300 58590
rect 880 58370 1300 58552
rect 58684 58370 59200 58590
rect 880 58280 59200 58370
rect 880 58272 59120 58280
rect 800 58000 59120 58272
rect 800 57600 59200 58000
rect 880 57510 59120 57600
rect 880 57320 1300 57510
rect 800 57290 1300 57320
rect 58684 57320 59120 57510
rect 58684 57290 59200 57320
rect 800 56920 59200 57290
rect 800 56648 59120 56920
rect 880 56640 59120 56648
rect 880 56430 59200 56640
rect 880 56368 1300 56430
rect 800 56210 1300 56368
rect 58684 56240 59200 56430
rect 58684 56210 59120 56240
rect 800 55960 59120 56210
rect 800 55560 59200 55960
rect 880 55350 59120 55560
rect 880 55280 1300 55350
rect 800 55130 1300 55280
rect 58684 55280 59120 55350
rect 58684 55130 59200 55280
rect 800 54744 59200 55130
rect 800 54608 59120 54744
rect 880 54464 59120 54608
rect 880 54328 59200 54464
rect 800 54270 59200 54328
rect 800 54050 1300 54270
rect 58684 54064 59200 54270
rect 58684 54050 59120 54064
rect 800 53784 59120 54050
rect 800 53656 59200 53784
rect 880 53384 59200 53656
rect 880 53376 59120 53384
rect 800 53190 59120 53376
rect 800 52970 1300 53190
rect 58684 53104 59120 53190
rect 58684 52970 59200 53104
rect 800 52704 59200 52970
rect 880 52424 59120 52704
rect 800 52110 59200 52424
rect 800 51890 1300 52110
rect 58684 52024 59200 52110
rect 58684 51890 59120 52024
rect 800 51744 59120 51890
rect 800 51616 59200 51744
rect 880 51344 59200 51616
rect 880 51336 59120 51344
rect 800 51064 59120 51336
rect 800 51030 59200 51064
rect 800 50810 1300 51030
rect 58684 50810 59200 51030
rect 800 50664 59200 50810
rect 880 50384 59120 50664
rect 800 49984 59200 50384
rect 800 49950 59120 49984
rect 800 49730 1300 49950
rect 58684 49730 59120 49950
rect 800 49712 59120 49730
rect 880 49704 59120 49712
rect 880 49432 59200 49704
rect 800 49168 59200 49432
rect 800 48888 59120 49168
rect 800 48870 59200 48888
rect 800 48760 1300 48870
rect 880 48650 1300 48760
rect 58684 48650 59200 48870
rect 880 48488 59200 48650
rect 880 48480 59120 48488
rect 800 48208 59120 48480
rect 800 47808 59200 48208
rect 880 47790 59120 47808
rect 880 47570 1300 47790
rect 58684 47570 59120 47790
rect 880 47528 59120 47570
rect 800 47128 59200 47528
rect 800 46848 59120 47128
rect 800 46720 59200 46848
rect 880 46710 59200 46720
rect 880 46490 1300 46710
rect 58684 46490 59200 46710
rect 880 46448 59200 46490
rect 880 46440 59120 46448
rect 800 46168 59120 46440
rect 800 45768 59200 46168
rect 880 45630 59120 45768
rect 880 45488 1300 45630
rect 800 45410 1300 45488
rect 58684 45488 59120 45630
rect 58684 45410 59200 45488
rect 800 45088 59200 45410
rect 800 44816 59120 45088
rect 880 44808 59120 44816
rect 880 44550 59200 44808
rect 880 44536 1300 44550
rect 800 44330 1300 44536
rect 58684 44408 59200 44550
rect 58684 44330 59120 44408
rect 800 44128 59120 44330
rect 800 43864 59200 44128
rect 880 43592 59200 43864
rect 880 43584 59120 43592
rect 800 43470 59120 43584
rect 800 43250 1300 43470
rect 58684 43312 59120 43470
rect 58684 43250 59200 43312
rect 800 42912 59200 43250
rect 800 42776 59120 42912
rect 880 42632 59120 42776
rect 880 42496 59200 42632
rect 800 42390 59200 42496
rect 800 42170 1300 42390
rect 58684 42232 59200 42390
rect 58684 42170 59120 42232
rect 800 41952 59120 42170
rect 800 41824 59200 41952
rect 880 41552 59200 41824
rect 880 41544 59120 41552
rect 800 41310 59120 41544
rect 800 41090 1300 41310
rect 58684 41272 59120 41310
rect 58684 41090 59200 41272
rect 800 40872 59200 41090
rect 880 40592 59120 40872
rect 800 40230 59200 40592
rect 800 40010 1300 40230
rect 58684 40192 59200 40230
rect 58684 40010 59120 40192
rect 800 39920 59120 40010
rect 880 39912 59120 39920
rect 880 39640 59200 39912
rect 800 39512 59200 39640
rect 800 39232 59120 39512
rect 800 39150 59200 39232
rect 800 38930 1300 39150
rect 58684 38930 59200 39150
rect 800 38832 59200 38930
rect 880 38552 59120 38832
rect 800 38070 59200 38552
rect 800 37880 1300 38070
rect 58684 38016 59200 38070
rect 880 37850 1300 37880
rect 58684 37850 59120 38016
rect 880 37736 59120 37850
rect 880 37600 59200 37736
rect 800 37336 59200 37600
rect 800 37056 59120 37336
rect 800 36990 59200 37056
rect 800 36928 1300 36990
rect 880 36770 1300 36928
rect 58684 36770 59200 36990
rect 880 36656 59200 36770
rect 880 36648 59120 36656
rect 800 36376 59120 36648
rect 800 35976 59200 36376
rect 880 35910 59120 35976
rect 880 35696 1300 35910
rect 800 35690 1300 35696
rect 58684 35696 59120 35910
rect 58684 35690 59200 35696
rect 800 35296 59200 35690
rect 800 35024 59120 35296
rect 880 35016 59120 35024
rect 880 34830 59200 35016
rect 880 34744 1300 34830
rect 800 34610 1300 34744
rect 58684 34616 59200 34830
rect 58684 34610 59120 34616
rect 800 34336 59120 34610
rect 800 33936 59200 34336
rect 880 33750 59120 33936
rect 880 33656 1300 33750
rect 800 33530 1300 33656
rect 58684 33656 59120 33750
rect 58684 33530 59200 33656
rect 800 33256 59200 33530
rect 800 32984 59120 33256
rect 880 32976 59120 32984
rect 880 32704 59200 32976
rect 800 32670 59200 32704
rect 800 32450 1300 32670
rect 58684 32450 59200 32670
rect 800 32440 59200 32450
rect 800 32160 59120 32440
rect 800 32032 59200 32160
rect 880 31760 59200 32032
rect 880 31752 59120 31760
rect 800 31590 59120 31752
rect 800 31370 1300 31590
rect 58684 31480 59120 31590
rect 58684 31370 59200 31480
rect 800 31080 59200 31370
rect 880 30800 59120 31080
rect 800 30510 59200 30800
rect 800 30290 1300 30510
rect 58684 30400 59200 30510
rect 58684 30290 59120 30400
rect 800 30120 59120 30290
rect 800 29992 59200 30120
rect 880 29720 59200 29992
rect 880 29712 59120 29720
rect 800 29440 59120 29712
rect 800 29430 59200 29440
rect 800 29210 1300 29430
rect 58684 29210 59200 29430
rect 800 29040 59200 29210
rect 880 28760 59120 29040
rect 800 28360 59200 28760
rect 800 28350 59120 28360
rect 800 28130 1300 28350
rect 58684 28130 59120 28350
rect 800 28088 59120 28130
rect 880 28080 59120 28088
rect 880 27808 59200 28080
rect 800 27544 59200 27808
rect 800 27270 59120 27544
rect 800 27136 1300 27270
rect 58684 27264 59120 27270
rect 880 27050 1300 27136
rect 58684 27050 59200 27264
rect 880 26864 59200 27050
rect 880 26856 59120 26864
rect 800 26584 59120 26856
rect 800 26190 59200 26584
rect 800 26048 1300 26190
rect 58684 26184 59200 26190
rect 880 25970 1300 26048
rect 58684 25970 59120 26184
rect 880 25904 59120 25970
rect 880 25768 59200 25904
rect 800 25504 59200 25768
rect 800 25224 59120 25504
rect 800 25110 59200 25224
rect 800 25096 1300 25110
rect 880 24890 1300 25096
rect 58684 24890 59200 25110
rect 880 24824 59200 24890
rect 880 24816 59120 24824
rect 800 24544 59120 24816
rect 800 24144 59200 24544
rect 880 24030 59120 24144
rect 880 23864 1300 24030
rect 800 23810 1300 23864
rect 58684 23864 59120 24030
rect 58684 23810 59200 23864
rect 800 23464 59200 23810
rect 800 23192 59120 23464
rect 880 23184 59120 23192
rect 880 22950 59200 23184
rect 880 22912 1300 22950
rect 800 22730 1300 22912
rect 58684 22784 59200 22950
rect 58684 22730 59120 22784
rect 800 22504 59120 22730
rect 800 22240 59200 22504
rect 880 21968 59200 22240
rect 880 21960 59120 21968
rect 800 21870 59120 21960
rect 800 21650 1300 21870
rect 58684 21688 59120 21870
rect 58684 21650 59200 21688
rect 800 21288 59200 21650
rect 800 21152 59120 21288
rect 880 21008 59120 21152
rect 880 20872 59200 21008
rect 800 20790 59200 20872
rect 800 20570 1300 20790
rect 58684 20608 59200 20790
rect 58684 20570 59120 20608
rect 800 20328 59120 20570
rect 800 20200 59200 20328
rect 880 19928 59200 20200
rect 880 19920 59120 19928
rect 800 19710 59120 19920
rect 800 19490 1300 19710
rect 58684 19648 59120 19710
rect 58684 19490 59200 19648
rect 800 19248 59200 19490
rect 880 18968 59120 19248
rect 800 18630 59200 18968
rect 800 18410 1300 18630
rect 58684 18568 59200 18630
rect 58684 18410 59120 18568
rect 800 18296 59120 18410
rect 880 18288 59120 18296
rect 880 18016 59200 18288
rect 800 17888 59200 18016
rect 800 17608 59120 17888
rect 800 17550 59200 17608
rect 800 17330 1300 17550
rect 58684 17330 59200 17550
rect 800 17208 59200 17330
rect 880 16928 59120 17208
rect 800 16470 59200 16928
rect 800 16256 1300 16470
rect 58684 16392 59200 16470
rect 880 16250 1300 16256
rect 58684 16250 59120 16392
rect 880 16112 59120 16250
rect 880 15976 59200 16112
rect 800 15712 59200 15976
rect 800 15432 59120 15712
rect 800 15390 59200 15432
rect 800 15304 1300 15390
rect 880 15170 1300 15304
rect 58684 15170 59200 15390
rect 880 15032 59200 15170
rect 880 15024 59120 15032
rect 800 14752 59120 15024
rect 800 14352 59200 14752
rect 880 14310 59120 14352
rect 880 14090 1300 14310
rect 58684 14090 59120 14310
rect 880 14072 59120 14090
rect 800 13672 59200 14072
rect 800 13392 59120 13672
rect 800 13264 59200 13392
rect 880 13230 59200 13264
rect 880 13010 1300 13230
rect 58684 13010 59200 13230
rect 880 12992 59200 13010
rect 880 12984 59120 12992
rect 800 12712 59120 12984
rect 800 12312 59200 12712
rect 880 12150 59120 12312
rect 880 12032 1300 12150
rect 800 11930 1300 12032
rect 58684 12032 59120 12150
rect 58684 11930 59200 12032
rect 800 11632 59200 11930
rect 800 11360 59120 11632
rect 880 11352 59120 11360
rect 880 11080 59200 11352
rect 800 11070 59200 11080
rect 800 10850 1300 11070
rect 58684 10850 59200 11070
rect 800 10816 59200 10850
rect 800 10536 59120 10816
rect 800 10408 59200 10536
rect 880 10136 59200 10408
rect 880 10128 59120 10136
rect 800 9990 59120 10128
rect 800 9770 1300 9990
rect 58684 9856 59120 9990
rect 58684 9770 59200 9856
rect 800 9456 59200 9770
rect 880 9176 59120 9456
rect 800 8910 59200 9176
rect 800 8690 1300 8910
rect 58684 8776 59200 8910
rect 58684 8690 59120 8776
rect 800 8496 59120 8690
rect 800 8368 59200 8496
rect 880 8096 59200 8368
rect 880 8088 59120 8096
rect 800 7830 59120 8088
rect 800 7610 1300 7830
rect 58684 7816 59120 7830
rect 58684 7610 59200 7816
rect 800 7416 59200 7610
rect 880 7136 59120 7416
rect 800 6750 59200 7136
rect 800 6530 1300 6750
rect 58684 6736 59200 6750
rect 58684 6530 59120 6736
rect 800 6464 59120 6530
rect 880 6456 59120 6464
rect 880 6184 59200 6456
rect 800 6056 59200 6184
rect 800 5776 59120 6056
rect 800 5670 59200 5776
rect 800 5512 1300 5670
rect 880 5450 1300 5512
rect 58684 5450 59200 5670
rect 880 5240 59200 5450
rect 880 5232 59120 5240
rect 800 4960 59120 5232
rect 800 4590 59200 4960
rect 800 4424 1300 4590
rect 58684 4560 59200 4590
rect 880 4370 1300 4424
rect 58684 4370 59120 4560
rect 880 4280 59120 4370
rect 880 4144 59200 4280
rect 800 3880 59200 4144
rect 800 3600 59120 3880
rect 800 3510 59200 3600
rect 800 3472 1300 3510
rect 880 3290 1300 3472
rect 58684 3290 59200 3510
rect 880 3200 59200 3290
rect 880 3192 59120 3200
rect 800 2920 59120 3192
rect 800 2520 59200 2920
rect 880 2430 59120 2520
rect 880 2240 1300 2430
rect 800 2210 1300 2240
rect 58684 2240 59120 2430
rect 58684 2210 59200 2240
rect 800 1840 59200 2210
rect 800 1568 59120 1840
rect 880 1560 59120 1568
rect 880 1350 59200 1560
rect 880 1288 1300 1350
rect 800 1130 1300 1288
rect 58684 1160 59200 1350
rect 58684 1130 59120 1160
rect 800 880 59120 1130
rect 800 616 59200 880
rect 880 480 59200 616
rect 880 336 59120 480
rect 800 307 59120 336
<< labels >>
rlabel metal3 s 0 5312 800 5432 6 cfg_colbits[0]
port 1 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 cfg_colbits[1]
port 2 nsew signal output
rlabel metal3 s 0 20000 800 20120 6 cfg_req_depth[0]
port 3 nsew signal output
rlabel metal3 s 0 20952 800 21072 6 cfg_req_depth[1]
port 4 nsew signal output
rlabel metal3 s 0 34824 800 34944 6 cfg_sdr_cas[0]
port 5 nsew signal output
rlabel metal3 s 0 35776 800 35896 6 cfg_sdr_cas[1]
port 6 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 cfg_sdr_cas[2]
port 7 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 cfg_sdr_en
port 8 nsew signal output
rlabel metal3 s 0 22040 800 22160 6 cfg_sdr_mode_reg[0]
port 9 nsew signal output
rlabel metal3 s 0 31832 800 31952 6 cfg_sdr_mode_reg[10]
port 10 nsew signal output
rlabel metal3 s 0 32784 800 32904 6 cfg_sdr_mode_reg[11]
port 11 nsew signal output
rlabel metal3 s 0 33736 800 33856 6 cfg_sdr_mode_reg[12]
port 12 nsew signal output
rlabel metal3 s 0 22992 800 23112 6 cfg_sdr_mode_reg[1]
port 13 nsew signal output
rlabel metal3 s 0 23944 800 24064 6 cfg_sdr_mode_reg[2]
port 14 nsew signal output
rlabel metal3 s 0 24896 800 25016 6 cfg_sdr_mode_reg[3]
port 15 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 cfg_sdr_mode_reg[4]
port 16 nsew signal output
rlabel metal3 s 0 26936 800 27056 6 cfg_sdr_mode_reg[5]
port 17 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 cfg_sdr_mode_reg[6]
port 18 nsew signal output
rlabel metal3 s 0 28840 800 28960 6 cfg_sdr_mode_reg[7]
port 19 nsew signal output
rlabel metal3 s 0 29792 800 29912 6 cfg_sdr_mode_reg[8]
port 20 nsew signal output
rlabel metal3 s 0 30880 800 31000 6 cfg_sdr_mode_reg[9]
port 21 nsew signal output
rlabel metal3 s 0 57400 800 57520 6 cfg_sdr_rfmax[0]
port 22 nsew signal output
rlabel metal3 s 0 58352 800 58472 6 cfg_sdr_rfmax[1]
port 23 nsew signal output
rlabel metal3 s 0 59304 800 59424 6 cfg_sdr_rfmax[2]
port 24 nsew signal output
rlabel metal3 s 0 45568 800 45688 6 cfg_sdr_rfsh[0]
port 25 nsew signal output
rlabel metal3 s 0 55360 800 55480 6 cfg_sdr_rfsh[10]
port 26 nsew signal output
rlabel metal3 s 0 56448 800 56568 6 cfg_sdr_rfsh[11]
port 27 nsew signal output
rlabel metal3 s 0 46520 800 46640 6 cfg_sdr_rfsh[1]
port 28 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 cfg_sdr_rfsh[2]
port 29 nsew signal output
rlabel metal3 s 0 48560 800 48680 6 cfg_sdr_rfsh[3]
port 30 nsew signal output
rlabel metal3 s 0 49512 800 49632 6 cfg_sdr_rfsh[4]
port 31 nsew signal output
rlabel metal3 s 0 50464 800 50584 6 cfg_sdr_rfsh[5]
port 32 nsew signal output
rlabel metal3 s 0 51416 800 51536 6 cfg_sdr_rfsh[6]
port 33 nsew signal output
rlabel metal3 s 0 52504 800 52624 6 cfg_sdr_rfsh[7]
port 34 nsew signal output
rlabel metal3 s 0 53456 800 53576 6 cfg_sdr_rfsh[8]
port 35 nsew signal output
rlabel metal3 s 0 54408 800 54528 6 cfg_sdr_rfsh[9]
port 36 nsew signal output
rlabel metal3 s 0 7216 800 7336 6 cfg_sdr_tras_d[0]
port 37 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 cfg_sdr_tras_d[1]
port 38 nsew signal output
rlabel metal3 s 0 9256 800 9376 6 cfg_sdr_tras_d[2]
port 39 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 cfg_sdr_tras_d[3]
port 40 nsew signal output
rlabel metal3 s 0 37680 800 37800 6 cfg_sdr_trcar_d[0]
port 41 nsew signal output
rlabel metal3 s 0 38632 800 38752 6 cfg_sdr_trcar_d[1]
port 42 nsew signal output
rlabel metal3 s 0 39720 800 39840 6 cfg_sdr_trcar_d[2]
port 43 nsew signal output
rlabel metal3 s 0 40672 800 40792 6 cfg_sdr_trcar_d[3]
port 44 nsew signal output
rlabel metal3 s 0 15104 800 15224 6 cfg_sdr_trcd_d[0]
port 45 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 cfg_sdr_trcd_d[1]
port 46 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 cfg_sdr_trcd_d[2]
port 47 nsew signal output
rlabel metal3 s 0 18096 800 18216 6 cfg_sdr_trcd_d[3]
port 48 nsew signal output
rlabel metal3 s 0 11160 800 11280 6 cfg_sdr_trp_d[0]
port 49 nsew signal output
rlabel metal3 s 0 12112 800 12232 6 cfg_sdr_trp_d[1]
port 50 nsew signal output
rlabel metal3 s 0 13064 800 13184 6 cfg_sdr_trp_d[2]
port 51 nsew signal output
rlabel metal3 s 0 14152 800 14272 6 cfg_sdr_trp_d[3]
port 52 nsew signal output
rlabel metal3 s 0 41624 800 41744 6 cfg_sdr_twr_d[0]
port 53 nsew signal output
rlabel metal3 s 0 42576 800 42696 6 cfg_sdr_twr_d[1]
port 54 nsew signal output
rlabel metal3 s 0 43664 800 43784 6 cfg_sdr_twr_d[2]
port 55 nsew signal output
rlabel metal3 s 0 44616 800 44736 6 cfg_sdr_twr_d[3]
port 56 nsew signal output
rlabel metal3 s 0 3272 800 3392 6 cfg_sdr_width[0]
port 57 nsew signal output
rlabel metal3 s 0 4224 800 4344 6 cfg_sdr_width[1]
port 58 nsew signal output
rlabel metal3 s 59200 1640 60000 1760 6 cpu_rst_n
port 59 nsew signal output
rlabel metal3 s 59200 3000 60000 3120 6 device_idcode[0]
port 60 nsew signal output
rlabel metal3 s 59200 9936 60000 10056 6 device_idcode[10]
port 61 nsew signal output
rlabel metal3 s 59200 10616 60000 10736 6 device_idcode[11]
port 62 nsew signal output
rlabel metal3 s 59200 11432 60000 11552 6 device_idcode[12]
port 63 nsew signal output
rlabel metal3 s 59200 12112 60000 12232 6 device_idcode[13]
port 64 nsew signal output
rlabel metal3 s 59200 12792 60000 12912 6 device_idcode[14]
port 65 nsew signal output
rlabel metal3 s 59200 13472 60000 13592 6 device_idcode[15]
port 66 nsew signal output
rlabel metal3 s 59200 14152 60000 14272 6 device_idcode[16]
port 67 nsew signal output
rlabel metal3 s 59200 14832 60000 14952 6 device_idcode[17]
port 68 nsew signal output
rlabel metal3 s 59200 15512 60000 15632 6 device_idcode[18]
port 69 nsew signal output
rlabel metal3 s 59200 16192 60000 16312 6 device_idcode[19]
port 70 nsew signal output
rlabel metal3 s 59200 3680 60000 3800 6 device_idcode[1]
port 71 nsew signal output
rlabel metal3 s 59200 17008 60000 17128 6 device_idcode[20]
port 72 nsew signal output
rlabel metal3 s 59200 17688 60000 17808 6 device_idcode[21]
port 73 nsew signal output
rlabel metal3 s 59200 18368 60000 18488 6 device_idcode[22]
port 74 nsew signal output
rlabel metal3 s 59200 19048 60000 19168 6 device_idcode[23]
port 75 nsew signal output
rlabel metal3 s 59200 19728 60000 19848 6 device_idcode[24]
port 76 nsew signal output
rlabel metal3 s 59200 20408 60000 20528 6 device_idcode[25]
port 77 nsew signal output
rlabel metal3 s 59200 21088 60000 21208 6 device_idcode[26]
port 78 nsew signal output
rlabel metal3 s 59200 21768 60000 21888 6 device_idcode[27]
port 79 nsew signal output
rlabel metal3 s 59200 22584 60000 22704 6 device_idcode[28]
port 80 nsew signal output
rlabel metal3 s 59200 23264 60000 23384 6 device_idcode[29]
port 81 nsew signal output
rlabel metal3 s 59200 4360 60000 4480 6 device_idcode[2]
port 82 nsew signal output
rlabel metal3 s 59200 23944 60000 24064 6 device_idcode[30]
port 83 nsew signal output
rlabel metal3 s 59200 24624 60000 24744 6 device_idcode[31]
port 84 nsew signal output
rlabel metal3 s 59200 5040 60000 5160 6 device_idcode[3]
port 85 nsew signal output
rlabel metal3 s 59200 5856 60000 5976 6 device_idcode[4]
port 86 nsew signal output
rlabel metal3 s 59200 6536 60000 6656 6 device_idcode[5]
port 87 nsew signal output
rlabel metal3 s 59200 7216 60000 7336 6 device_idcode[6]
port 88 nsew signal output
rlabel metal3 s 59200 7896 60000 8016 6 device_idcode[7]
port 89 nsew signal output
rlabel metal3 s 59200 8576 60000 8696 6 device_idcode[8]
port 90 nsew signal output
rlabel metal3 s 59200 9256 60000 9376 6 device_idcode[9]
port 91 nsew signal output
rlabel metal3 s 59200 25304 60000 25424 6 fuse_mhartid[0]
port 92 nsew signal output
rlabel metal3 s 59200 32240 60000 32360 6 fuse_mhartid[10]
port 93 nsew signal output
rlabel metal3 s 59200 33056 60000 33176 6 fuse_mhartid[11]
port 94 nsew signal output
rlabel metal3 s 59200 33736 60000 33856 6 fuse_mhartid[12]
port 95 nsew signal output
rlabel metal3 s 59200 34416 60000 34536 6 fuse_mhartid[13]
port 96 nsew signal output
rlabel metal3 s 59200 35096 60000 35216 6 fuse_mhartid[14]
port 97 nsew signal output
rlabel metal3 s 59200 35776 60000 35896 6 fuse_mhartid[15]
port 98 nsew signal output
rlabel metal3 s 59200 36456 60000 36576 6 fuse_mhartid[16]
port 99 nsew signal output
rlabel metal3 s 59200 37136 60000 37256 6 fuse_mhartid[17]
port 100 nsew signal output
rlabel metal3 s 59200 37816 60000 37936 6 fuse_mhartid[18]
port 101 nsew signal output
rlabel metal3 s 59200 38632 60000 38752 6 fuse_mhartid[19]
port 102 nsew signal output
rlabel metal3 s 59200 25984 60000 26104 6 fuse_mhartid[1]
port 103 nsew signal output
rlabel metal3 s 59200 39312 60000 39432 6 fuse_mhartid[20]
port 104 nsew signal output
rlabel metal3 s 59200 39992 60000 40112 6 fuse_mhartid[21]
port 105 nsew signal output
rlabel metal3 s 59200 40672 60000 40792 6 fuse_mhartid[22]
port 106 nsew signal output
rlabel metal3 s 59200 41352 60000 41472 6 fuse_mhartid[23]
port 107 nsew signal output
rlabel metal3 s 59200 42032 60000 42152 6 fuse_mhartid[24]
port 108 nsew signal output
rlabel metal3 s 59200 42712 60000 42832 6 fuse_mhartid[25]
port 109 nsew signal output
rlabel metal3 s 59200 43392 60000 43512 6 fuse_mhartid[26]
port 110 nsew signal output
rlabel metal3 s 59200 44208 60000 44328 6 fuse_mhartid[27]
port 111 nsew signal output
rlabel metal3 s 59200 44888 60000 45008 6 fuse_mhartid[28]
port 112 nsew signal output
rlabel metal3 s 59200 45568 60000 45688 6 fuse_mhartid[29]
port 113 nsew signal output
rlabel metal3 s 59200 26664 60000 26784 6 fuse_mhartid[2]
port 114 nsew signal output
rlabel metal3 s 59200 46248 60000 46368 6 fuse_mhartid[30]
port 115 nsew signal output
rlabel metal3 s 59200 46928 60000 47048 6 fuse_mhartid[31]
port 116 nsew signal output
rlabel metal3 s 59200 27344 60000 27464 6 fuse_mhartid[3]
port 117 nsew signal output
rlabel metal3 s 59200 28160 60000 28280 6 fuse_mhartid[4]
port 118 nsew signal output
rlabel metal3 s 59200 28840 60000 28960 6 fuse_mhartid[5]
port 119 nsew signal output
rlabel metal3 s 59200 29520 60000 29640 6 fuse_mhartid[6]
port 120 nsew signal output
rlabel metal3 s 59200 30200 60000 30320 6 fuse_mhartid[7]
port 121 nsew signal output
rlabel metal3 s 59200 30880 60000 31000 6 fuse_mhartid[8]
port 122 nsew signal output
rlabel metal3 s 59200 31560 60000 31680 6 fuse_mhartid[9]
port 123 nsew signal output
rlabel metal3 s 59200 47608 60000 47728 6 irq_lines[0]
port 124 nsew signal output
rlabel metal3 s 59200 54544 60000 54664 6 irq_lines[10]
port 125 nsew signal output
rlabel metal3 s 59200 55360 60000 55480 6 irq_lines[11]
port 126 nsew signal output
rlabel metal3 s 59200 56040 60000 56160 6 irq_lines[12]
port 127 nsew signal output
rlabel metal3 s 59200 56720 60000 56840 6 irq_lines[13]
port 128 nsew signal output
rlabel metal3 s 59200 57400 60000 57520 6 irq_lines[14]
port 129 nsew signal output
rlabel metal3 s 59200 58080 60000 58200 6 irq_lines[15]
port 130 nsew signal output
rlabel metal3 s 59200 48288 60000 48408 6 irq_lines[1]
port 131 nsew signal output
rlabel metal3 s 59200 48968 60000 49088 6 irq_lines[2]
port 132 nsew signal output
rlabel metal3 s 59200 49784 60000 49904 6 irq_lines[3]
port 133 nsew signal output
rlabel metal3 s 59200 50464 60000 50584 6 irq_lines[4]
port 134 nsew signal output
rlabel metal3 s 59200 51144 60000 51264 6 irq_lines[5]
port 135 nsew signal output
rlabel metal3 s 59200 51824 60000 51944 6 irq_lines[6]
port 136 nsew signal output
rlabel metal3 s 59200 52504 60000 52624 6 irq_lines[7]
port 137 nsew signal output
rlabel metal3 s 59200 53184 60000 53304 6 irq_lines[8]
port 138 nsew signal output
rlabel metal3 s 59200 53864 60000 53984 6 irq_lines[9]
port 139 nsew signal output
rlabel metal3 s 59200 280 60000 400 6 mclk
port 140 nsew signal input
rlabel metal2 s 58714 59200 58770 60000 6 reg_ack
port 141 nsew signal output
rlabel metal2 s 1950 59200 2006 60000 6 reg_addr[0]
port 142 nsew signal input
rlabel metal2 s 2686 59200 2742 60000 6 reg_addr[1]
port 143 nsew signal input
rlabel metal2 s 3514 59200 3570 60000 6 reg_addr[2]
port 144 nsew signal input
rlabel metal2 s 4250 59200 4306 60000 6 reg_addr[3]
port 145 nsew signal input
rlabel metal2 s 5078 59200 5134 60000 6 reg_be[0]
port 146 nsew signal input
rlabel metal2 s 5906 59200 5962 60000 6 reg_be[1]
port 147 nsew signal input
rlabel metal2 s 6642 59200 6698 60000 6 reg_be[2]
port 148 nsew signal input
rlabel metal2 s 7470 59200 7526 60000 6 reg_be[3]
port 149 nsew signal input
rlabel metal2 s 386 59200 442 60000 6 reg_cs
port 150 nsew signal input
rlabel metal2 s 33506 59200 33562 60000 6 reg_rdata[0]
port 151 nsew signal output
rlabel metal2 s 41418 59200 41474 60000 6 reg_rdata[10]
port 152 nsew signal output
rlabel metal2 s 42154 59200 42210 60000 6 reg_rdata[11]
port 153 nsew signal output
rlabel metal2 s 42982 59200 43038 60000 6 reg_rdata[12]
port 154 nsew signal output
rlabel metal2 s 43718 59200 43774 60000 6 reg_rdata[13]
port 155 nsew signal output
rlabel metal2 s 44546 59200 44602 60000 6 reg_rdata[14]
port 156 nsew signal output
rlabel metal2 s 45374 59200 45430 60000 6 reg_rdata[15]
port 157 nsew signal output
rlabel metal2 s 46110 59200 46166 60000 6 reg_rdata[16]
port 158 nsew signal output
rlabel metal2 s 46938 59200 46994 60000 6 reg_rdata[17]
port 159 nsew signal output
rlabel metal2 s 47674 59200 47730 60000 6 reg_rdata[18]
port 160 nsew signal output
rlabel metal2 s 48502 59200 48558 60000 6 reg_rdata[19]
port 161 nsew signal output
rlabel metal2 s 34242 59200 34298 60000 6 reg_rdata[1]
port 162 nsew signal output
rlabel metal2 s 49238 59200 49294 60000 6 reg_rdata[20]
port 163 nsew signal output
rlabel metal2 s 50066 59200 50122 60000 6 reg_rdata[21]
port 164 nsew signal output
rlabel metal2 s 50894 59200 50950 60000 6 reg_rdata[22]
port 165 nsew signal output
rlabel metal2 s 51630 59200 51686 60000 6 reg_rdata[23]
port 166 nsew signal output
rlabel metal2 s 52458 59200 52514 60000 6 reg_rdata[24]
port 167 nsew signal output
rlabel metal2 s 53194 59200 53250 60000 6 reg_rdata[25]
port 168 nsew signal output
rlabel metal2 s 54022 59200 54078 60000 6 reg_rdata[26]
port 169 nsew signal output
rlabel metal2 s 54758 59200 54814 60000 6 reg_rdata[27]
port 170 nsew signal output
rlabel metal2 s 55586 59200 55642 60000 6 reg_rdata[28]
port 171 nsew signal output
rlabel metal2 s 56414 59200 56470 60000 6 reg_rdata[29]
port 172 nsew signal output
rlabel metal2 s 35070 59200 35126 60000 6 reg_rdata[2]
port 173 nsew signal output
rlabel metal2 s 57150 59200 57206 60000 6 reg_rdata[30]
port 174 nsew signal output
rlabel metal2 s 57978 59200 58034 60000 6 reg_rdata[31]
port 175 nsew signal output
rlabel metal2 s 35898 59200 35954 60000 6 reg_rdata[3]
port 176 nsew signal output
rlabel metal2 s 36634 59200 36690 60000 6 reg_rdata[4]
port 177 nsew signal output
rlabel metal2 s 37462 59200 37518 60000 6 reg_rdata[5]
port 178 nsew signal output
rlabel metal2 s 38198 59200 38254 60000 6 reg_rdata[6]
port 179 nsew signal output
rlabel metal2 s 39026 59200 39082 60000 6 reg_rdata[7]
port 180 nsew signal output
rlabel metal2 s 39762 59200 39818 60000 6 reg_rdata[8]
port 181 nsew signal output
rlabel metal2 s 40590 59200 40646 60000 6 reg_rdata[9]
port 182 nsew signal output
rlabel metal2 s 8206 59200 8262 60000 6 reg_wdata[0]
port 183 nsew signal input
rlabel metal2 s 16118 59200 16174 60000 6 reg_wdata[10]
port 184 nsew signal input
rlabel metal2 s 16946 59200 17002 60000 6 reg_wdata[11]
port 185 nsew signal input
rlabel metal2 s 17682 59200 17738 60000 6 reg_wdata[12]
port 186 nsew signal input
rlabel metal2 s 18510 59200 18566 60000 6 reg_wdata[13]
port 187 nsew signal input
rlabel metal2 s 19246 59200 19302 60000 6 reg_wdata[14]
port 188 nsew signal input
rlabel metal2 s 20074 59200 20130 60000 6 reg_wdata[15]
port 189 nsew signal input
rlabel metal2 s 20902 59200 20958 60000 6 reg_wdata[16]
port 190 nsew signal input
rlabel metal2 s 21638 59200 21694 60000 6 reg_wdata[17]
port 191 nsew signal input
rlabel metal2 s 22466 59200 22522 60000 6 reg_wdata[18]
port 192 nsew signal input
rlabel metal2 s 23202 59200 23258 60000 6 reg_wdata[19]
port 193 nsew signal input
rlabel metal2 s 9034 59200 9090 60000 6 reg_wdata[1]
port 194 nsew signal input
rlabel metal2 s 24030 59200 24086 60000 6 reg_wdata[20]
port 195 nsew signal input
rlabel metal2 s 24766 59200 24822 60000 6 reg_wdata[21]
port 196 nsew signal input
rlabel metal2 s 25594 59200 25650 60000 6 reg_wdata[22]
port 197 nsew signal input
rlabel metal2 s 26422 59200 26478 60000 6 reg_wdata[23]
port 198 nsew signal input
rlabel metal2 s 27158 59200 27214 60000 6 reg_wdata[24]
port 199 nsew signal input
rlabel metal2 s 27986 59200 28042 60000 6 reg_wdata[25]
port 200 nsew signal input
rlabel metal2 s 28722 59200 28778 60000 6 reg_wdata[26]
port 201 nsew signal input
rlabel metal2 s 29550 59200 29606 60000 6 reg_wdata[27]
port 202 nsew signal input
rlabel metal2 s 30378 59200 30434 60000 6 reg_wdata[28]
port 203 nsew signal input
rlabel metal2 s 31114 59200 31170 60000 6 reg_wdata[29]
port 204 nsew signal input
rlabel metal2 s 9770 59200 9826 60000 6 reg_wdata[2]
port 205 nsew signal input
rlabel metal2 s 31942 59200 31998 60000 6 reg_wdata[30]
port 206 nsew signal input
rlabel metal2 s 32678 59200 32734 60000 6 reg_wdata[31]
port 207 nsew signal input
rlabel metal2 s 10598 59200 10654 60000 6 reg_wdata[3]
port 208 nsew signal input
rlabel metal2 s 11426 59200 11482 60000 6 reg_wdata[4]
port 209 nsew signal input
rlabel metal2 s 12162 59200 12218 60000 6 reg_wdata[5]
port 210 nsew signal input
rlabel metal2 s 12990 59200 13046 60000 6 reg_wdata[6]
port 211 nsew signal input
rlabel metal2 s 13726 59200 13782 60000 6 reg_wdata[7]
port 212 nsew signal input
rlabel metal2 s 14554 59200 14610 60000 6 reg_wdata[8]
port 213 nsew signal input
rlabel metal2 s 15382 59200 15438 60000 6 reg_wdata[9]
port 214 nsew signal input
rlabel metal2 s 1122 59200 1178 60000 6 reg_wr
port 215 nsew signal input
rlabel metal3 s 59200 960 60000 1080 6 reset_n
port 216 nsew signal input
rlabel metal3 s 0 2320 800 2440 6 sdr_init_done
port 217 nsew signal input
rlabel metal3 s 0 416 800 536 6 sdram_clk
port 218 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 sdram_rst_n
port 219 nsew signal output
rlabel metal3 s 59200 58760 60000 58880 6 soft_irq
port 220 nsew signal output
rlabel metal3 s 59200 2320 60000 2440 6 spi_rst_n
port 221 nsew signal output
rlabel metal2 s 30010 0 30066 800 6 user_irq[0]
port 222 nsew signal output
rlabel metal3 s 59200 59440 60000 59560 6 user_irq[1]
port 223 nsew signal output
rlabel metal2 s 59542 59200 59598 60000 6 user_irq[2]
port 224 nsew signal output
rlabel metal2 s 51350 1040 51410 58800 6 VPWR
port 225 nsew power bidirectional
rlabel metal2 s 35350 1040 35410 58800 6 VPWR
port 226 nsew power bidirectional
rlabel metal2 s 19350 1040 19410 58800 6 VPWR
port 227 nsew power bidirectional
rlabel metal2 s 3350 1040 3410 58800 6 VPWR
port 228 nsew power bidirectional
rlabel metal3 s 1380 57370 58604 57430 6 VPWR
port 229 nsew power bidirectional
rlabel metal3 s 1380 55210 58604 55270 6 VPWR
port 230 nsew power bidirectional
rlabel metal3 s 1380 53050 58604 53110 6 VPWR
port 231 nsew power bidirectional
rlabel metal3 s 1380 50890 58604 50950 6 VPWR
port 232 nsew power bidirectional
rlabel metal3 s 1380 48730 58604 48790 6 VPWR
port 233 nsew power bidirectional
rlabel metal3 s 1380 46570 58604 46630 6 VPWR
port 234 nsew power bidirectional
rlabel metal3 s 1380 44410 58604 44470 6 VPWR
port 235 nsew power bidirectional
rlabel metal3 s 1380 42250 58604 42310 6 VPWR
port 236 nsew power bidirectional
rlabel metal3 s 1380 40090 58604 40150 6 VPWR
port 237 nsew power bidirectional
rlabel metal3 s 1380 37930 58604 37990 6 VPWR
port 238 nsew power bidirectional
rlabel metal3 s 1380 35770 58604 35830 6 VPWR
port 239 nsew power bidirectional
rlabel metal3 s 1380 33610 58604 33670 6 VPWR
port 240 nsew power bidirectional
rlabel metal3 s 1380 31450 58604 31510 6 VPWR
port 241 nsew power bidirectional
rlabel metal3 s 1380 29290 58604 29350 6 VPWR
port 242 nsew power bidirectional
rlabel metal3 s 1380 27130 58604 27190 6 VPWR
port 243 nsew power bidirectional
rlabel metal3 s 1380 24970 58604 25030 6 VPWR
port 244 nsew power bidirectional
rlabel metal3 s 1380 22810 58604 22870 6 VPWR
port 245 nsew power bidirectional
rlabel metal3 s 1380 20650 58604 20710 6 VPWR
port 246 nsew power bidirectional
rlabel metal3 s 1380 18490 58604 18550 6 VPWR
port 247 nsew power bidirectional
rlabel metal3 s 1380 16330 58604 16390 6 VPWR
port 248 nsew power bidirectional
rlabel metal3 s 1380 14170 58604 14230 6 VPWR
port 249 nsew power bidirectional
rlabel metal3 s 1380 12010 58604 12070 6 VPWR
port 250 nsew power bidirectional
rlabel metal3 s 1380 9850 58604 9910 6 VPWR
port 251 nsew power bidirectional
rlabel metal3 s 1380 7690 58604 7750 6 VPWR
port 252 nsew power bidirectional
rlabel metal3 s 1380 5530 58604 5590 6 VPWR
port 253 nsew power bidirectional
rlabel metal3 s 1380 3370 58604 3430 6 VPWR
port 254 nsew power bidirectional
rlabel metal3 s 1380 1210 58604 1270 6 VPWR
port 255 nsew power bidirectional
rlabel metal2 s 43350 1040 43410 58800 6 VGND
port 256 nsew ground bidirectional
rlabel metal2 s 27350 1040 27410 58800 6 VGND
port 257 nsew ground bidirectional
rlabel metal2 s 11350 1040 11410 58800 6 VGND
port 258 nsew ground bidirectional
rlabel metal3 s 1380 58450 58604 58510 6 VGND
port 259 nsew ground bidirectional
rlabel metal3 s 1380 56290 58604 56350 6 VGND
port 260 nsew ground bidirectional
rlabel metal3 s 1380 54130 58604 54190 6 VGND
port 261 nsew ground bidirectional
rlabel metal3 s 1380 51970 58604 52030 6 VGND
port 262 nsew ground bidirectional
rlabel metal3 s 1380 49810 58604 49870 6 VGND
port 263 nsew ground bidirectional
rlabel metal3 s 1380 47650 58604 47710 6 VGND
port 264 nsew ground bidirectional
rlabel metal3 s 1380 45490 58604 45550 6 VGND
port 265 nsew ground bidirectional
rlabel metal3 s 1380 43330 58604 43390 6 VGND
port 266 nsew ground bidirectional
rlabel metal3 s 1380 41170 58604 41230 6 VGND
port 267 nsew ground bidirectional
rlabel metal3 s 1380 39010 58604 39070 6 VGND
port 268 nsew ground bidirectional
rlabel metal3 s 1380 36850 58604 36910 6 VGND
port 269 nsew ground bidirectional
rlabel metal3 s 1380 34690 58604 34750 6 VGND
port 270 nsew ground bidirectional
rlabel metal3 s 1380 32530 58604 32590 6 VGND
port 271 nsew ground bidirectional
rlabel metal3 s 1380 30370 58604 30430 6 VGND
port 272 nsew ground bidirectional
rlabel metal3 s 1380 28210 58604 28270 6 VGND
port 273 nsew ground bidirectional
rlabel metal3 s 1380 26050 58604 26110 6 VGND
port 274 nsew ground bidirectional
rlabel metal3 s 1380 23890 58604 23950 6 VGND
port 275 nsew ground bidirectional
rlabel metal3 s 1380 21730 58604 21790 6 VGND
port 276 nsew ground bidirectional
rlabel metal3 s 1380 19570 58604 19630 6 VGND
port 277 nsew ground bidirectional
rlabel metal3 s 1380 17410 58604 17470 6 VGND
port 278 nsew ground bidirectional
rlabel metal3 s 1380 15250 58604 15310 6 VGND
port 279 nsew ground bidirectional
rlabel metal3 s 1380 13090 58604 13150 6 VGND
port 280 nsew ground bidirectional
rlabel metal3 s 1380 10930 58604 10990 6 VGND
port 281 nsew ground bidirectional
rlabel metal3 s 1380 8770 58604 8830 6 VGND
port 282 nsew ground bidirectional
rlabel metal3 s 1380 6610 58604 6670 6 VGND
port 283 nsew ground bidirectional
rlabel metal3 s 1380 4450 58604 4510 6 VGND
port 284 nsew ground bidirectional
rlabel metal3 s 1380 2290 58604 2350 6 VGND
port 285 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 60000 60000
string LEFview TRUE
string GDS_FILE /project/openlane/glbl_cfg/runs/glbl_cfg/results/magic/glbl_cfg.gds
string GDS_END 7483434
string GDS_START 184298
<< end >>

