magic
tech sky130A
magscale 1 2
timestamp 1623948498
<< obsli1 >>
rect 1104 2159 198812 57681
<< obsm1 >>
rect 934 2048 199074 57996
<< metal2 >>
rect 938 59200 994 60000
rect 2778 59200 2834 60000
rect 4710 59200 4766 60000
rect 6550 59200 6606 60000
rect 8482 59200 8538 60000
rect 10322 59200 10378 60000
rect 12254 59200 12310 60000
rect 14094 59200 14150 60000
rect 16026 59200 16082 60000
rect 17866 59200 17922 60000
rect 19798 59200 19854 60000
rect 21638 59200 21694 60000
rect 23570 59200 23626 60000
rect 25410 59200 25466 60000
rect 27342 59200 27398 60000
rect 29182 59200 29238 60000
rect 31114 59200 31170 60000
rect 32954 59200 33010 60000
rect 34886 59200 34942 60000
rect 36726 59200 36782 60000
rect 38658 59200 38714 60000
rect 40498 59200 40554 60000
rect 42430 59200 42486 60000
rect 44270 59200 44326 60000
rect 46202 59200 46258 60000
rect 48042 59200 48098 60000
rect 49974 59200 50030 60000
rect 51814 59200 51870 60000
rect 53746 59200 53802 60000
rect 55586 59200 55642 60000
rect 57518 59200 57574 60000
rect 59358 59200 59414 60000
rect 61290 59200 61346 60000
rect 63130 59200 63186 60000
rect 65062 59200 65118 60000
rect 66902 59200 66958 60000
rect 68834 59200 68890 60000
rect 70674 59200 70730 60000
rect 72606 59200 72662 60000
rect 74446 59200 74502 60000
rect 76378 59200 76434 60000
rect 78218 59200 78274 60000
rect 80150 59200 80206 60000
rect 81990 59200 82046 60000
rect 83922 59200 83978 60000
rect 85762 59200 85818 60000
rect 87694 59200 87750 60000
rect 89534 59200 89590 60000
rect 91466 59200 91522 60000
rect 93306 59200 93362 60000
rect 95238 59200 95294 60000
rect 97078 59200 97134 60000
rect 99010 59200 99066 60000
rect 100942 59200 100998 60000
rect 102782 59200 102838 60000
rect 104714 59200 104770 60000
rect 106554 59200 106610 60000
rect 108486 59200 108542 60000
rect 110326 59200 110382 60000
rect 112258 59200 112314 60000
rect 114098 59200 114154 60000
rect 116030 59200 116086 60000
rect 117870 59200 117926 60000
rect 119802 59200 119858 60000
rect 121642 59200 121698 60000
rect 123574 59200 123630 60000
rect 125414 59200 125470 60000
rect 127346 59200 127402 60000
rect 129186 59200 129242 60000
rect 131118 59200 131174 60000
rect 132958 59200 133014 60000
rect 134890 59200 134946 60000
rect 136730 59200 136786 60000
rect 138662 59200 138718 60000
rect 140502 59200 140558 60000
rect 142434 59200 142490 60000
rect 144274 59200 144330 60000
rect 146206 59200 146262 60000
rect 148046 59200 148102 60000
rect 149978 59200 150034 60000
rect 151818 59200 151874 60000
rect 153750 59200 153806 60000
rect 155590 59200 155646 60000
rect 157522 59200 157578 60000
rect 159362 59200 159418 60000
rect 161294 59200 161350 60000
rect 163134 59200 163190 60000
rect 165066 59200 165122 60000
rect 166906 59200 166962 60000
rect 168838 59200 168894 60000
rect 170678 59200 170734 60000
rect 172610 59200 172666 60000
rect 174450 59200 174506 60000
rect 176382 59200 176438 60000
rect 178222 59200 178278 60000
rect 180154 59200 180210 60000
rect 181994 59200 182050 60000
rect 183926 59200 183982 60000
rect 185766 59200 185822 60000
rect 187698 59200 187754 60000
rect 189538 59200 189594 60000
rect 191470 59200 191526 60000
rect 193310 59200 193366 60000
rect 195242 59200 195298 60000
rect 197082 59200 197138 60000
rect 199014 59200 199070 60000
rect 2502 0 2558 800
rect 7562 0 7618 800
rect 12714 0 12770 800
rect 17866 0 17922 800
rect 22926 0 22982 800
rect 28078 0 28134 800
rect 33230 0 33286 800
rect 38382 0 38438 800
rect 43442 0 43498 800
rect 48594 0 48650 800
rect 53746 0 53802 800
rect 58898 0 58954 800
rect 63958 0 64014 800
rect 69110 0 69166 800
rect 74262 0 74318 800
rect 79414 0 79470 800
rect 84474 0 84530 800
rect 89626 0 89682 800
rect 94778 0 94834 800
rect 99930 0 99986 800
rect 104990 0 105046 800
rect 110142 0 110198 800
rect 115294 0 115350 800
rect 120446 0 120502 800
rect 125506 0 125562 800
rect 130658 0 130714 800
rect 135810 0 135866 800
rect 140962 0 141018 800
rect 146022 0 146078 800
rect 151174 0 151230 800
rect 156326 0 156382 800
rect 161478 0 161534 800
rect 166538 0 166594 800
rect 171690 0 171746 800
rect 176842 0 176898 800
rect 181994 0 182050 800
rect 187054 0 187110 800
rect 192206 0 192262 800
rect 197358 0 197414 800
<< obsm2 >>
rect 1050 59144 2722 59401
rect 2890 59144 4654 59401
rect 4822 59144 6494 59401
rect 6662 59144 8426 59401
rect 8594 59144 10266 59401
rect 10434 59144 12198 59401
rect 12366 59144 14038 59401
rect 14206 59144 15970 59401
rect 16138 59144 17810 59401
rect 17978 59144 19742 59401
rect 19910 59144 21582 59401
rect 21750 59144 23514 59401
rect 23682 59144 25354 59401
rect 25522 59144 27286 59401
rect 27454 59144 29126 59401
rect 29294 59144 31058 59401
rect 31226 59144 32898 59401
rect 33066 59144 34830 59401
rect 34998 59144 36670 59401
rect 36838 59144 38602 59401
rect 38770 59144 40442 59401
rect 40610 59144 42374 59401
rect 42542 59144 44214 59401
rect 44382 59144 46146 59401
rect 46314 59144 47986 59401
rect 48154 59144 49918 59401
rect 50086 59144 51758 59401
rect 51926 59144 53690 59401
rect 53858 59144 55530 59401
rect 55698 59144 57462 59401
rect 57630 59144 59302 59401
rect 59470 59144 61234 59401
rect 61402 59144 63074 59401
rect 63242 59144 65006 59401
rect 65174 59144 66846 59401
rect 67014 59144 68778 59401
rect 68946 59144 70618 59401
rect 70786 59144 72550 59401
rect 72718 59144 74390 59401
rect 74558 59144 76322 59401
rect 76490 59144 78162 59401
rect 78330 59144 80094 59401
rect 80262 59144 81934 59401
rect 82102 59144 83866 59401
rect 84034 59144 85706 59401
rect 85874 59144 87638 59401
rect 87806 59144 89478 59401
rect 89646 59144 91410 59401
rect 91578 59144 93250 59401
rect 93418 59144 95182 59401
rect 95350 59144 97022 59401
rect 97190 59144 98954 59401
rect 99122 59144 100886 59401
rect 101054 59144 102726 59401
rect 102894 59144 104658 59401
rect 104826 59144 106498 59401
rect 106666 59144 108430 59401
rect 108598 59144 110270 59401
rect 110438 59144 112202 59401
rect 112370 59144 114042 59401
rect 114210 59144 115974 59401
rect 116142 59144 117814 59401
rect 117982 59144 119746 59401
rect 119914 59144 121586 59401
rect 121754 59144 123518 59401
rect 123686 59144 125358 59401
rect 125526 59144 127290 59401
rect 127458 59144 129130 59401
rect 129298 59144 131062 59401
rect 131230 59144 132902 59401
rect 133070 59144 134834 59401
rect 135002 59144 136674 59401
rect 136842 59144 138606 59401
rect 138774 59144 140446 59401
rect 140614 59144 142378 59401
rect 142546 59144 144218 59401
rect 144386 59144 146150 59401
rect 146318 59144 147990 59401
rect 148158 59144 149922 59401
rect 150090 59144 151762 59401
rect 151930 59144 153694 59401
rect 153862 59144 155534 59401
rect 155702 59144 157466 59401
rect 157634 59144 159306 59401
rect 159474 59144 161238 59401
rect 161406 59144 163078 59401
rect 163246 59144 165010 59401
rect 165178 59144 166850 59401
rect 167018 59144 168782 59401
rect 168950 59144 170622 59401
rect 170790 59144 172554 59401
rect 172722 59144 174394 59401
rect 174562 59144 176326 59401
rect 176494 59144 178166 59401
rect 178334 59144 180098 59401
rect 180266 59144 181938 59401
rect 182106 59144 183870 59401
rect 184038 59144 185710 59401
rect 185878 59144 187642 59401
rect 187810 59144 189482 59401
rect 189650 59144 191414 59401
rect 191582 59144 193254 59401
rect 193422 59144 195186 59401
rect 195354 59144 197026 59401
rect 197194 59144 198958 59401
rect 940 856 199068 59144
rect 940 439 2446 856
rect 2614 439 7506 856
rect 7674 439 12658 856
rect 12826 439 17810 856
rect 17978 439 22870 856
rect 23038 439 28022 856
rect 28190 439 33174 856
rect 33342 439 38326 856
rect 38494 439 43386 856
rect 43554 439 48538 856
rect 48706 439 53690 856
rect 53858 439 58842 856
rect 59010 439 63902 856
rect 64070 439 69054 856
rect 69222 439 74206 856
rect 74374 439 79358 856
rect 79526 439 84418 856
rect 84586 439 89570 856
rect 89738 439 94722 856
rect 94890 439 99874 856
rect 100042 439 104934 856
rect 105102 439 110086 856
rect 110254 439 115238 856
rect 115406 439 120390 856
rect 120558 439 125450 856
rect 125618 439 130602 856
rect 130770 439 135754 856
rect 135922 439 140906 856
rect 141074 439 145966 856
rect 146134 439 151118 856
rect 151286 439 156270 856
rect 156438 439 161422 856
rect 161590 439 166482 856
rect 166650 439 171634 856
rect 171802 439 176786 856
rect 176954 439 181938 856
rect 182106 439 186998 856
rect 187166 439 192150 856
rect 192318 439 197302 856
rect 197470 439 199068 856
<< metal3 >>
rect 199200 59304 200000 59424
rect 199200 58352 200000 58472
rect 199200 57400 200000 57520
rect 199200 56448 200000 56568
rect 199200 55360 200000 55480
rect 199200 54408 200000 54528
rect 199200 53456 200000 53576
rect 199200 52504 200000 52624
rect 199200 51416 200000 51536
rect 199200 50464 200000 50584
rect 0 49920 800 50040
rect 199200 49512 200000 49632
rect 199200 48560 200000 48680
rect 199200 47608 200000 47728
rect 199200 46520 200000 46640
rect 199200 45568 200000 45688
rect 199200 44616 200000 44736
rect 199200 43664 200000 43784
rect 199200 42576 200000 42696
rect 199200 41624 200000 41744
rect 199200 40672 200000 40792
rect 199200 39720 200000 39840
rect 199200 38632 200000 38752
rect 199200 37680 200000 37800
rect 199200 36728 200000 36848
rect 199200 35776 200000 35896
rect 199200 34824 200000 34944
rect 199200 33736 200000 33856
rect 199200 32784 200000 32904
rect 199200 31832 200000 31952
rect 199200 30880 200000 31000
rect 0 29928 800 30048
rect 199200 29792 200000 29912
rect 199200 28840 200000 28960
rect 199200 27888 200000 28008
rect 199200 26936 200000 27056
rect 199200 25848 200000 25968
rect 199200 24896 200000 25016
rect 199200 23944 200000 24064
rect 199200 22992 200000 23112
rect 199200 22040 200000 22160
rect 199200 20952 200000 21072
rect 199200 20000 200000 20120
rect 199200 19048 200000 19168
rect 199200 18096 200000 18216
rect 199200 17008 200000 17128
rect 199200 16056 200000 16176
rect 199200 15104 200000 15224
rect 199200 14152 200000 14272
rect 199200 13064 200000 13184
rect 199200 12112 200000 12232
rect 199200 11160 200000 11280
rect 199200 10208 200000 10328
rect 0 9936 800 10056
rect 199200 9256 200000 9376
rect 199200 8168 200000 8288
rect 199200 7216 200000 7336
rect 199200 6264 200000 6384
rect 199200 5312 200000 5432
rect 199200 4224 200000 4344
rect 199200 3272 200000 3392
rect 199200 2320 200000 2440
rect 199200 1368 200000 1488
rect 199200 416 200000 536
<< obsm3 >>
rect 800 59224 199120 59397
rect 800 58552 199200 59224
rect 800 58272 199120 58552
rect 800 57600 199200 58272
rect 800 57320 199120 57600
rect 800 56648 199200 57320
rect 800 56368 199120 56648
rect 800 55560 199200 56368
rect 800 55280 199120 55560
rect 800 54608 199200 55280
rect 800 54328 199120 54608
rect 800 53656 199200 54328
rect 800 53376 199120 53656
rect 800 52704 199200 53376
rect 800 52424 199120 52704
rect 800 51616 199200 52424
rect 800 51336 199120 51616
rect 800 50664 199200 51336
rect 800 50384 199120 50664
rect 800 50120 199200 50384
rect 880 49840 199200 50120
rect 800 49712 199200 49840
rect 800 49432 199120 49712
rect 800 48760 199200 49432
rect 800 48480 199120 48760
rect 800 47808 199200 48480
rect 800 47528 199120 47808
rect 800 46720 199200 47528
rect 800 46440 199120 46720
rect 800 45768 199200 46440
rect 800 45488 199120 45768
rect 800 44816 199200 45488
rect 800 44536 199120 44816
rect 800 43864 199200 44536
rect 800 43584 199120 43864
rect 800 42776 199200 43584
rect 800 42496 199120 42776
rect 800 41824 199200 42496
rect 800 41544 199120 41824
rect 800 40872 199200 41544
rect 800 40592 199120 40872
rect 800 39920 199200 40592
rect 800 39640 199120 39920
rect 800 38832 199200 39640
rect 800 38552 199120 38832
rect 800 37880 199200 38552
rect 800 37600 199120 37880
rect 800 36928 199200 37600
rect 800 36648 199120 36928
rect 800 35976 199200 36648
rect 800 35696 199120 35976
rect 800 35024 199200 35696
rect 800 34744 199120 35024
rect 800 33936 199200 34744
rect 800 33656 199120 33936
rect 800 32984 199200 33656
rect 800 32704 199120 32984
rect 800 32032 199200 32704
rect 800 31752 199120 32032
rect 800 31080 199200 31752
rect 800 30800 199120 31080
rect 800 30128 199200 30800
rect 880 29992 199200 30128
rect 880 29848 199120 29992
rect 800 29712 199120 29848
rect 800 29040 199200 29712
rect 800 28760 199120 29040
rect 800 28088 199200 28760
rect 800 27808 199120 28088
rect 800 27136 199200 27808
rect 800 26856 199120 27136
rect 800 26048 199200 26856
rect 800 25768 199120 26048
rect 800 25096 199200 25768
rect 800 24816 199120 25096
rect 800 24144 199200 24816
rect 800 23864 199120 24144
rect 800 23192 199200 23864
rect 800 22912 199120 23192
rect 800 22240 199200 22912
rect 800 21960 199120 22240
rect 800 21152 199200 21960
rect 800 20872 199120 21152
rect 800 20200 199200 20872
rect 800 19920 199120 20200
rect 800 19248 199200 19920
rect 800 18968 199120 19248
rect 800 18296 199200 18968
rect 800 18016 199120 18296
rect 800 17208 199200 18016
rect 800 16928 199120 17208
rect 800 16256 199200 16928
rect 800 15976 199120 16256
rect 800 15304 199200 15976
rect 800 15024 199120 15304
rect 800 14352 199200 15024
rect 800 14072 199120 14352
rect 800 13264 199200 14072
rect 800 12984 199120 13264
rect 800 12312 199200 12984
rect 800 12032 199120 12312
rect 800 11360 199200 12032
rect 800 11080 199120 11360
rect 800 10408 199200 11080
rect 800 10136 199120 10408
rect 880 10128 199120 10136
rect 880 9856 199200 10128
rect 800 9456 199200 9856
rect 800 9176 199120 9456
rect 800 8368 199200 9176
rect 800 8088 199120 8368
rect 800 7416 199200 8088
rect 800 7136 199120 7416
rect 800 6464 199200 7136
rect 800 6184 199120 6464
rect 800 5512 199200 6184
rect 800 5232 199120 5512
rect 800 4424 199200 5232
rect 800 4144 199120 4424
rect 800 3472 199200 4144
rect 800 3192 199120 3472
rect 800 2520 199200 3192
rect 800 2240 199120 2520
rect 800 1568 199200 2240
rect 800 1288 199120 1568
rect 800 616 199200 1288
rect 800 443 199120 616
<< metal4 >>
rect 4208 2128 4528 57712
rect 19568 2128 19888 57712
rect 34928 2128 35248 57712
rect 50288 2128 50608 57712
rect 65648 2128 65968 57712
rect 81008 2128 81328 57712
rect 96368 2128 96688 57712
rect 111728 2128 112048 57712
rect 127088 2128 127408 57712
rect 142448 2128 142768 57712
rect 157808 2128 158128 57712
rect 173168 2128 173488 57712
rect 188528 2128 188848 57712
<< labels >>
rlabel metal3 s 199200 3272 200000 3392 6 cfg_colbits[0]
port 1 nsew signal input
rlabel metal3 s 199200 4224 200000 4344 6 cfg_colbits[1]
port 2 nsew signal input
rlabel metal3 s 199200 18096 200000 18216 6 cfg_req_depth[0]
port 3 nsew signal input
rlabel metal3 s 199200 19048 200000 19168 6 cfg_req_depth[1]
port 4 nsew signal input
rlabel metal3 s 199200 32784 200000 32904 6 cfg_sdr_cas[0]
port 5 nsew signal input
rlabel metal3 s 199200 33736 200000 33856 6 cfg_sdr_cas[1]
port 6 nsew signal input
rlabel metal3 s 199200 34824 200000 34944 6 cfg_sdr_cas[2]
port 7 nsew signal input
rlabel metal3 s 199200 17008 200000 17128 6 cfg_sdr_en
port 8 nsew signal input
rlabel metal3 s 199200 20000 200000 20120 6 cfg_sdr_mode_reg[0]
port 9 nsew signal input
rlabel metal3 s 199200 29792 200000 29912 6 cfg_sdr_mode_reg[10]
port 10 nsew signal input
rlabel metal3 s 199200 30880 200000 31000 6 cfg_sdr_mode_reg[11]
port 11 nsew signal input
rlabel metal3 s 199200 31832 200000 31952 6 cfg_sdr_mode_reg[12]
port 12 nsew signal input
rlabel metal3 s 199200 20952 200000 21072 6 cfg_sdr_mode_reg[1]
port 13 nsew signal input
rlabel metal3 s 199200 22040 200000 22160 6 cfg_sdr_mode_reg[2]
port 14 nsew signal input
rlabel metal3 s 199200 22992 200000 23112 6 cfg_sdr_mode_reg[3]
port 15 nsew signal input
rlabel metal3 s 199200 23944 200000 24064 6 cfg_sdr_mode_reg[4]
port 16 nsew signal input
rlabel metal3 s 199200 24896 200000 25016 6 cfg_sdr_mode_reg[5]
port 17 nsew signal input
rlabel metal3 s 199200 25848 200000 25968 6 cfg_sdr_mode_reg[6]
port 18 nsew signal input
rlabel metal3 s 199200 26936 200000 27056 6 cfg_sdr_mode_reg[7]
port 19 nsew signal input
rlabel metal3 s 199200 27888 200000 28008 6 cfg_sdr_mode_reg[8]
port 20 nsew signal input
rlabel metal3 s 199200 28840 200000 28960 6 cfg_sdr_mode_reg[9]
port 21 nsew signal input
rlabel metal3 s 199200 55360 200000 55480 6 cfg_sdr_rfmax[0]
port 22 nsew signal input
rlabel metal3 s 199200 56448 200000 56568 6 cfg_sdr_rfmax[1]
port 23 nsew signal input
rlabel metal3 s 199200 57400 200000 57520 6 cfg_sdr_rfmax[2]
port 24 nsew signal input
rlabel metal3 s 199200 43664 200000 43784 6 cfg_sdr_rfsh[0]
port 25 nsew signal input
rlabel metal3 s 199200 53456 200000 53576 6 cfg_sdr_rfsh[10]
port 26 nsew signal input
rlabel metal3 s 199200 54408 200000 54528 6 cfg_sdr_rfsh[11]
port 27 nsew signal input
rlabel metal3 s 199200 44616 200000 44736 6 cfg_sdr_rfsh[1]
port 28 nsew signal input
rlabel metal3 s 199200 45568 200000 45688 6 cfg_sdr_rfsh[2]
port 29 nsew signal input
rlabel metal3 s 199200 46520 200000 46640 6 cfg_sdr_rfsh[3]
port 30 nsew signal input
rlabel metal3 s 199200 47608 200000 47728 6 cfg_sdr_rfsh[4]
port 31 nsew signal input
rlabel metal3 s 199200 48560 200000 48680 6 cfg_sdr_rfsh[5]
port 32 nsew signal input
rlabel metal3 s 199200 49512 200000 49632 6 cfg_sdr_rfsh[6]
port 33 nsew signal input
rlabel metal3 s 199200 50464 200000 50584 6 cfg_sdr_rfsh[7]
port 34 nsew signal input
rlabel metal3 s 199200 51416 200000 51536 6 cfg_sdr_rfsh[8]
port 35 nsew signal input
rlabel metal3 s 199200 52504 200000 52624 6 cfg_sdr_rfsh[9]
port 36 nsew signal input
rlabel metal3 s 199200 5312 200000 5432 6 cfg_sdr_tras_d[0]
port 37 nsew signal input
rlabel metal3 s 199200 6264 200000 6384 6 cfg_sdr_tras_d[1]
port 38 nsew signal input
rlabel metal3 s 199200 7216 200000 7336 6 cfg_sdr_tras_d[2]
port 39 nsew signal input
rlabel metal3 s 199200 8168 200000 8288 6 cfg_sdr_tras_d[3]
port 40 nsew signal input
rlabel metal3 s 199200 35776 200000 35896 6 cfg_sdr_trcar_d[0]
port 41 nsew signal input
rlabel metal3 s 199200 36728 200000 36848 6 cfg_sdr_trcar_d[1]
port 42 nsew signal input
rlabel metal3 s 199200 37680 200000 37800 6 cfg_sdr_trcar_d[2]
port 43 nsew signal input
rlabel metal3 s 199200 38632 200000 38752 6 cfg_sdr_trcar_d[3]
port 44 nsew signal input
rlabel metal3 s 199200 13064 200000 13184 6 cfg_sdr_trcd_d[0]
port 45 nsew signal input
rlabel metal3 s 199200 14152 200000 14272 6 cfg_sdr_trcd_d[1]
port 46 nsew signal input
rlabel metal3 s 199200 15104 200000 15224 6 cfg_sdr_trcd_d[2]
port 47 nsew signal input
rlabel metal3 s 199200 16056 200000 16176 6 cfg_sdr_trcd_d[3]
port 48 nsew signal input
rlabel metal3 s 199200 9256 200000 9376 6 cfg_sdr_trp_d[0]
port 49 nsew signal input
rlabel metal3 s 199200 10208 200000 10328 6 cfg_sdr_trp_d[1]
port 50 nsew signal input
rlabel metal3 s 199200 11160 200000 11280 6 cfg_sdr_trp_d[2]
port 51 nsew signal input
rlabel metal3 s 199200 12112 200000 12232 6 cfg_sdr_trp_d[3]
port 52 nsew signal input
rlabel metal3 s 199200 39720 200000 39840 6 cfg_sdr_twr_d[0]
port 53 nsew signal input
rlabel metal3 s 199200 40672 200000 40792 6 cfg_sdr_twr_d[1]
port 54 nsew signal input
rlabel metal3 s 199200 41624 200000 41744 6 cfg_sdr_twr_d[2]
port 55 nsew signal input
rlabel metal3 s 199200 42576 200000 42696 6 cfg_sdr_twr_d[3]
port 56 nsew signal input
rlabel metal3 s 199200 1368 200000 1488 6 cfg_sdr_width[0]
port 57 nsew signal input
rlabel metal3 s 199200 2320 200000 2440 6 cfg_sdr_width[1]
port 58 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 pad_sdr_din[0]
port 59 nsew signal input
rlabel metal2 s 84474 0 84530 800 6 pad_sdr_din[1]
port 60 nsew signal input
rlabel metal2 s 89626 0 89682 800 6 pad_sdr_din[2]
port 61 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 pad_sdr_din[3]
port 62 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 pad_sdr_din[4]
port 63 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 pad_sdr_din[5]
port 64 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 pad_sdr_din[6]
port 65 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 pad_sdr_din[7]
port 66 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 sdr_addr[0]
port 67 nsew signal output
rlabel metal2 s 53746 0 53802 800 6 sdr_addr[10]
port 68 nsew signal output
rlabel metal2 s 58898 0 58954 800 6 sdr_addr[11]
port 69 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 sdr_addr[12]
port 70 nsew signal output
rlabel metal2 s 7562 0 7618 800 6 sdr_addr[1]
port 71 nsew signal output
rlabel metal2 s 12714 0 12770 800 6 sdr_addr[2]
port 72 nsew signal output
rlabel metal2 s 17866 0 17922 800 6 sdr_addr[3]
port 73 nsew signal output
rlabel metal2 s 22926 0 22982 800 6 sdr_addr[4]
port 74 nsew signal output
rlabel metal2 s 28078 0 28134 800 6 sdr_addr[5]
port 75 nsew signal output
rlabel metal2 s 33230 0 33286 800 6 sdr_addr[6]
port 76 nsew signal output
rlabel metal2 s 38382 0 38438 800 6 sdr_addr[7]
port 77 nsew signal output
rlabel metal2 s 43442 0 43498 800 6 sdr_addr[8]
port 78 nsew signal output
rlabel metal2 s 48594 0 48650 800 6 sdr_addr[9]
port 79 nsew signal output
rlabel metal2 s 69110 0 69166 800 6 sdr_ba[0]
port 80 nsew signal output
rlabel metal2 s 74262 0 74318 800 6 sdr_ba[1]
port 81 nsew signal output
rlabel metal2 s 161478 0 161534 800 6 sdr_cas_n
port 82 nsew signal output
rlabel metal3 s 199200 58352 200000 58472 6 sdr_cke
port 83 nsew signal output
rlabel metal3 s 0 9936 800 10056 6 sdr_cs_n
port 84 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 sdr_den_n
port 85 nsew signal output
rlabel metal2 s 120446 0 120502 800 6 sdr_dout[0]
port 86 nsew signal output
rlabel metal2 s 125506 0 125562 800 6 sdr_dout[1]
port 87 nsew signal output
rlabel metal2 s 130658 0 130714 800 6 sdr_dout[2]
port 88 nsew signal output
rlabel metal2 s 135810 0 135866 800 6 sdr_dout[3]
port 89 nsew signal output
rlabel metal2 s 140962 0 141018 800 6 sdr_dout[4]
port 90 nsew signal output
rlabel metal2 s 146022 0 146078 800 6 sdr_dout[5]
port 91 nsew signal output
rlabel metal2 s 151174 0 151230 800 6 sdr_dout[6]
port 92 nsew signal output
rlabel metal2 s 156326 0 156382 800 6 sdr_dout[7]
port 93 nsew signal output
rlabel metal2 s 166538 0 166594 800 6 sdr_dqm
port 94 nsew signal output
rlabel metal2 s 171690 0 171746 800 6 sdr_init_done
port 95 nsew signal output
rlabel metal2 s 195242 59200 195298 60000 6 sdr_ras_n
port 96 nsew signal output
rlabel metal2 s 197082 59200 197138 60000 6 sdr_we_n
port 97 nsew signal output
rlabel metal2 s 176842 0 176898 800 6 sdram_clk
port 98 nsew signal input
rlabel metal2 s 199014 59200 199070 60000 6 sdram_pad_clk
port 99 nsew signal input
rlabel metal3 s 199200 416 200000 536 6 sdram_resetn
port 100 nsew signal input
rlabel metal3 s 0 49920 800 50040 6 wb_ack_o
port 101 nsew signal output
rlabel metal2 s 938 59200 994 60000 6 wb_addr_i[0]
port 102 nsew signal input
rlabel metal2 s 19798 59200 19854 60000 6 wb_addr_i[10]
port 103 nsew signal input
rlabel metal2 s 21638 59200 21694 60000 6 wb_addr_i[11]
port 104 nsew signal input
rlabel metal2 s 23570 59200 23626 60000 6 wb_addr_i[12]
port 105 nsew signal input
rlabel metal2 s 25410 59200 25466 60000 6 wb_addr_i[13]
port 106 nsew signal input
rlabel metal2 s 27342 59200 27398 60000 6 wb_addr_i[14]
port 107 nsew signal input
rlabel metal2 s 29182 59200 29238 60000 6 wb_addr_i[15]
port 108 nsew signal input
rlabel metal2 s 31114 59200 31170 60000 6 wb_addr_i[16]
port 109 nsew signal input
rlabel metal2 s 32954 59200 33010 60000 6 wb_addr_i[17]
port 110 nsew signal input
rlabel metal2 s 34886 59200 34942 60000 6 wb_addr_i[18]
port 111 nsew signal input
rlabel metal2 s 36726 59200 36782 60000 6 wb_addr_i[19]
port 112 nsew signal input
rlabel metal2 s 2778 59200 2834 60000 6 wb_addr_i[1]
port 113 nsew signal input
rlabel metal2 s 38658 59200 38714 60000 6 wb_addr_i[20]
port 114 nsew signal input
rlabel metal2 s 40498 59200 40554 60000 6 wb_addr_i[21]
port 115 nsew signal input
rlabel metal2 s 42430 59200 42486 60000 6 wb_addr_i[22]
port 116 nsew signal input
rlabel metal2 s 44270 59200 44326 60000 6 wb_addr_i[23]
port 117 nsew signal input
rlabel metal2 s 46202 59200 46258 60000 6 wb_addr_i[24]
port 118 nsew signal input
rlabel metal2 s 48042 59200 48098 60000 6 wb_addr_i[25]
port 119 nsew signal input
rlabel metal2 s 49974 59200 50030 60000 6 wb_addr_i[26]
port 120 nsew signal input
rlabel metal2 s 51814 59200 51870 60000 6 wb_addr_i[27]
port 121 nsew signal input
rlabel metal2 s 53746 59200 53802 60000 6 wb_addr_i[28]
port 122 nsew signal input
rlabel metal2 s 55586 59200 55642 60000 6 wb_addr_i[29]
port 123 nsew signal input
rlabel metal2 s 4710 59200 4766 60000 6 wb_addr_i[2]
port 124 nsew signal input
rlabel metal2 s 57518 59200 57574 60000 6 wb_addr_i[30]
port 125 nsew signal input
rlabel metal2 s 59358 59200 59414 60000 6 wb_addr_i[31]
port 126 nsew signal input
rlabel metal2 s 6550 59200 6606 60000 6 wb_addr_i[3]
port 127 nsew signal input
rlabel metal2 s 8482 59200 8538 60000 6 wb_addr_i[4]
port 128 nsew signal input
rlabel metal2 s 10322 59200 10378 60000 6 wb_addr_i[5]
port 129 nsew signal input
rlabel metal2 s 12254 59200 12310 60000 6 wb_addr_i[6]
port 130 nsew signal input
rlabel metal2 s 14094 59200 14150 60000 6 wb_addr_i[7]
port 131 nsew signal input
rlabel metal2 s 16026 59200 16082 60000 6 wb_addr_i[8]
port 132 nsew signal input
rlabel metal2 s 17866 59200 17922 60000 6 wb_addr_i[9]
port 133 nsew signal input
rlabel metal2 s 181994 0 182050 800 6 wb_clk_i
port 134 nsew signal input
rlabel metal2 s 189538 59200 189594 60000 6 wb_cti_i[0]
port 135 nsew signal input
rlabel metal2 s 191470 59200 191526 60000 6 wb_cti_i[1]
port 136 nsew signal input
rlabel metal2 s 193310 59200 193366 60000 6 wb_cti_i[2]
port 137 nsew signal input
rlabel metal3 s 199200 59304 200000 59424 6 wb_cyc_i
port 138 nsew signal input
rlabel metal2 s 68834 59200 68890 60000 6 wb_dat_i[0]
port 139 nsew signal input
rlabel metal2 s 87694 59200 87750 60000 6 wb_dat_i[10]
port 140 nsew signal input
rlabel metal2 s 89534 59200 89590 60000 6 wb_dat_i[11]
port 141 nsew signal input
rlabel metal2 s 91466 59200 91522 60000 6 wb_dat_i[12]
port 142 nsew signal input
rlabel metal2 s 93306 59200 93362 60000 6 wb_dat_i[13]
port 143 nsew signal input
rlabel metal2 s 95238 59200 95294 60000 6 wb_dat_i[14]
port 144 nsew signal input
rlabel metal2 s 97078 59200 97134 60000 6 wb_dat_i[15]
port 145 nsew signal input
rlabel metal2 s 99010 59200 99066 60000 6 wb_dat_i[16]
port 146 nsew signal input
rlabel metal2 s 100942 59200 100998 60000 6 wb_dat_i[17]
port 147 nsew signal input
rlabel metal2 s 102782 59200 102838 60000 6 wb_dat_i[18]
port 148 nsew signal input
rlabel metal2 s 104714 59200 104770 60000 6 wb_dat_i[19]
port 149 nsew signal input
rlabel metal2 s 70674 59200 70730 60000 6 wb_dat_i[1]
port 150 nsew signal input
rlabel metal2 s 106554 59200 106610 60000 6 wb_dat_i[20]
port 151 nsew signal input
rlabel metal2 s 108486 59200 108542 60000 6 wb_dat_i[21]
port 152 nsew signal input
rlabel metal2 s 110326 59200 110382 60000 6 wb_dat_i[22]
port 153 nsew signal input
rlabel metal2 s 112258 59200 112314 60000 6 wb_dat_i[23]
port 154 nsew signal input
rlabel metal2 s 114098 59200 114154 60000 6 wb_dat_i[24]
port 155 nsew signal input
rlabel metal2 s 116030 59200 116086 60000 6 wb_dat_i[25]
port 156 nsew signal input
rlabel metal2 s 117870 59200 117926 60000 6 wb_dat_i[26]
port 157 nsew signal input
rlabel metal2 s 119802 59200 119858 60000 6 wb_dat_i[27]
port 158 nsew signal input
rlabel metal2 s 121642 59200 121698 60000 6 wb_dat_i[28]
port 159 nsew signal input
rlabel metal2 s 123574 59200 123630 60000 6 wb_dat_i[29]
port 160 nsew signal input
rlabel metal2 s 72606 59200 72662 60000 6 wb_dat_i[2]
port 161 nsew signal input
rlabel metal2 s 125414 59200 125470 60000 6 wb_dat_i[30]
port 162 nsew signal input
rlabel metal2 s 127346 59200 127402 60000 6 wb_dat_i[31]
port 163 nsew signal input
rlabel metal2 s 74446 59200 74502 60000 6 wb_dat_i[3]
port 164 nsew signal input
rlabel metal2 s 76378 59200 76434 60000 6 wb_dat_i[4]
port 165 nsew signal input
rlabel metal2 s 78218 59200 78274 60000 6 wb_dat_i[5]
port 166 nsew signal input
rlabel metal2 s 80150 59200 80206 60000 6 wb_dat_i[6]
port 167 nsew signal input
rlabel metal2 s 81990 59200 82046 60000 6 wb_dat_i[7]
port 168 nsew signal input
rlabel metal2 s 83922 59200 83978 60000 6 wb_dat_i[8]
port 169 nsew signal input
rlabel metal2 s 85762 59200 85818 60000 6 wb_dat_i[9]
port 170 nsew signal input
rlabel metal2 s 129186 59200 129242 60000 6 wb_dat_o[0]
port 171 nsew signal output
rlabel metal2 s 148046 59200 148102 60000 6 wb_dat_o[10]
port 172 nsew signal output
rlabel metal2 s 149978 59200 150034 60000 6 wb_dat_o[11]
port 173 nsew signal output
rlabel metal2 s 151818 59200 151874 60000 6 wb_dat_o[12]
port 174 nsew signal output
rlabel metal2 s 153750 59200 153806 60000 6 wb_dat_o[13]
port 175 nsew signal output
rlabel metal2 s 155590 59200 155646 60000 6 wb_dat_o[14]
port 176 nsew signal output
rlabel metal2 s 157522 59200 157578 60000 6 wb_dat_o[15]
port 177 nsew signal output
rlabel metal2 s 159362 59200 159418 60000 6 wb_dat_o[16]
port 178 nsew signal output
rlabel metal2 s 161294 59200 161350 60000 6 wb_dat_o[17]
port 179 nsew signal output
rlabel metal2 s 163134 59200 163190 60000 6 wb_dat_o[18]
port 180 nsew signal output
rlabel metal2 s 165066 59200 165122 60000 6 wb_dat_o[19]
port 181 nsew signal output
rlabel metal2 s 131118 59200 131174 60000 6 wb_dat_o[1]
port 182 nsew signal output
rlabel metal2 s 166906 59200 166962 60000 6 wb_dat_o[20]
port 183 nsew signal output
rlabel metal2 s 168838 59200 168894 60000 6 wb_dat_o[21]
port 184 nsew signal output
rlabel metal2 s 170678 59200 170734 60000 6 wb_dat_o[22]
port 185 nsew signal output
rlabel metal2 s 172610 59200 172666 60000 6 wb_dat_o[23]
port 186 nsew signal output
rlabel metal2 s 174450 59200 174506 60000 6 wb_dat_o[24]
port 187 nsew signal output
rlabel metal2 s 176382 59200 176438 60000 6 wb_dat_o[25]
port 188 nsew signal output
rlabel metal2 s 178222 59200 178278 60000 6 wb_dat_o[26]
port 189 nsew signal output
rlabel metal2 s 180154 59200 180210 60000 6 wb_dat_o[27]
port 190 nsew signal output
rlabel metal2 s 181994 59200 182050 60000 6 wb_dat_o[28]
port 191 nsew signal output
rlabel metal2 s 183926 59200 183982 60000 6 wb_dat_o[29]
port 192 nsew signal output
rlabel metal2 s 132958 59200 133014 60000 6 wb_dat_o[2]
port 193 nsew signal output
rlabel metal2 s 185766 59200 185822 60000 6 wb_dat_o[30]
port 194 nsew signal output
rlabel metal2 s 187698 59200 187754 60000 6 wb_dat_o[31]
port 195 nsew signal output
rlabel metal2 s 134890 59200 134946 60000 6 wb_dat_o[3]
port 196 nsew signal output
rlabel metal2 s 136730 59200 136786 60000 6 wb_dat_o[4]
port 197 nsew signal output
rlabel metal2 s 138662 59200 138718 60000 6 wb_dat_o[5]
port 198 nsew signal output
rlabel metal2 s 140502 59200 140558 60000 6 wb_dat_o[6]
port 199 nsew signal output
rlabel metal2 s 142434 59200 142490 60000 6 wb_dat_o[7]
port 200 nsew signal output
rlabel metal2 s 144274 59200 144330 60000 6 wb_dat_o[8]
port 201 nsew signal output
rlabel metal2 s 146206 59200 146262 60000 6 wb_dat_o[9]
port 202 nsew signal output
rlabel metal2 s 187054 0 187110 800 6 wb_rst_i
port 203 nsew signal input
rlabel metal2 s 61290 59200 61346 60000 6 wb_sel_i[0]
port 204 nsew signal input
rlabel metal2 s 63130 59200 63186 60000 6 wb_sel_i[1]
port 205 nsew signal input
rlabel metal2 s 65062 59200 65118 60000 6 wb_sel_i[2]
port 206 nsew signal input
rlabel metal2 s 66902 59200 66958 60000 6 wb_sel_i[3]
port 207 nsew signal input
rlabel metal2 s 192206 0 192262 800 6 wb_stb_i
port 208 nsew signal input
rlabel metal2 s 197358 0 197414 800 6 wb_we_i
port 209 nsew signal input
rlabel metal4 s 188528 2128 188848 57712 6 VPWR
port 210 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 57712 6 VPWR
port 211 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 57712 6 VPWR
port 212 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 57712 6 VPWR
port 213 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 57712 6 VPWR
port 214 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 57712 6 VPWR
port 215 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 57712 6 VPWR
port 216 nsew power bidirectional
rlabel metal4 s 173168 2128 173488 57712 6 VGND
port 217 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 57712 6 VGND
port 218 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 57712 6 VGND
port 219 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 57712 6 VGND
port 220 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 57712 6 VGND
port 221 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 57712 6 VGND
port 222 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 200000 60000
string LEFview TRUE
string GDS_FILE /project/openlane/sdram/runs/sdram/results/magic/sdrc_top.gds
string GDS_END 17975034
string GDS_START 271150
<< end >>

