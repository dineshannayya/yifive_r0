module user_project_wrapper (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    vccd1,
    vssd1,
    vccd2,
    vssd2,
    vdda1,
    vssa1,
    vdda2,
    vssa2,
    analog_io,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input vccd1;
 input vssd1;
 input vccd2;
 input vssd2;
 input vdda1;
 input vssa1;
 input vdda2;
 input vssa2;
 inout [28:0] analog_io;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 sky130_fd_sc_hd__inv_4 _008_ (.A(wb_rst_i),
    .Y(\u_core.wb_rst_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _009_ (.A(\u_core.spi_en_tx ),
    .Y(io_oeb[35]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _010_ (.HI(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _011_ (.HI(io_oeb[37]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _012_ (.HI(_000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _013_ (.LO(_001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _014_ (.LO(_002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _015_ (.LO(la_data_out[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _016_ (.LO(la_data_out[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _017_ (.LO(la_data_out[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _018_ (.LO(la_data_out[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _019_ (.LO(la_data_out[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _020_ (.LO(la_data_out[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _021_ (.LO(la_data_out[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _022_ (.LO(la_data_out[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _023_ (.LO(la_data_out[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _024_ (.LO(la_data_out[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _025_ (.LO(la_data_out[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _026_ (.LO(la_data_out[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _027_ (.LO(la_data_out[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _028_ (.LO(la_data_out[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _029_ (.LO(la_data_out[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _030_ (.LO(la_data_out[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _031_ (.LO(la_data_out[16]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _032_ (.LO(la_data_out[17]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _033_ (.LO(la_data_out[18]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _034_ (.LO(la_data_out[19]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _035_ (.LO(la_data_out[20]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _036_ (.LO(la_data_out[21]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _037_ (.LO(la_data_out[22]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _038_ (.LO(la_data_out[23]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _039_ (.LO(la_data_out[24]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _040_ (.LO(la_data_out[25]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _041_ (.LO(la_data_out[26]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _042_ (.LO(la_data_out[27]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _043_ (.LO(la_data_out[28]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _044_ (.LO(la_data_out[29]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _045_ (.LO(la_data_out[30]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _046_ (.LO(la_data_out[31]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _047_ (.LO(la_data_out[32]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _048_ (.LO(la_data_out[33]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _049_ (.LO(la_data_out[34]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _050_ (.LO(la_data_out[35]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _051_ (.LO(la_data_out[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _052_ (.LO(la_data_out[37]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _053_ (.LO(la_data_out[38]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _054_ (.LO(la_data_out[39]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _055_ (.LO(la_data_out[40]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _056_ (.LO(la_data_out[41]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _057_ (.LO(la_data_out[42]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _058_ (.LO(la_data_out[43]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _059_ (.LO(la_data_out[44]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _060_ (.LO(la_data_out[45]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _061_ (.LO(la_data_out[46]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _062_ (.LO(la_data_out[47]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _063_ (.LO(la_data_out[48]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _064_ (.LO(la_data_out[49]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _065_ (.LO(la_data_out[50]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _066_ (.LO(la_data_out[51]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _067_ (.LO(la_data_out[52]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _068_ (.LO(la_data_out[53]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _069_ (.LO(la_data_out[54]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _070_ (.LO(la_data_out[55]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _071_ (.LO(la_data_out[56]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _072_ (.LO(la_data_out[57]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _073_ (.LO(la_data_out[58]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _074_ (.LO(la_data_out[59]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _075_ (.LO(la_data_out[60]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _076_ (.LO(la_data_out[61]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _077_ (.LO(la_data_out[62]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _078_ (.LO(la_data_out[63]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _079_ (.LO(la_data_out[64]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _080_ (.LO(la_data_out[65]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _081_ (.LO(la_data_out[66]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _082_ (.LO(la_data_out[67]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _083_ (.LO(la_data_out[68]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _084_ (.LO(la_data_out[69]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _085_ (.LO(la_data_out[70]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _086_ (.LO(la_data_out[71]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _087_ (.LO(la_data_out[72]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _088_ (.LO(la_data_out[73]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _089_ (.LO(la_data_out[74]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _090_ (.LO(la_data_out[75]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _091_ (.LO(la_data_out[76]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _092_ (.LO(la_data_out[77]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _093_ (.LO(la_data_out[78]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _094_ (.LO(la_data_out[79]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _095_ (.LO(la_data_out[80]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _096_ (.LO(la_data_out[81]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _097_ (.LO(la_data_out[82]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _098_ (.LO(la_data_out[83]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _099_ (.LO(la_data_out[84]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _100_ (.LO(la_data_out[85]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _101_ (.LO(la_data_out[86]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _102_ (.LO(la_data_out[87]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _103_ (.LO(la_data_out[88]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _104_ (.LO(la_data_out[89]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _105_ (.LO(la_data_out[90]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _106_ (.LO(la_data_out[91]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _107_ (.LO(la_data_out[92]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _108_ (.LO(la_data_out[93]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _109_ (.LO(la_data_out[94]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _110_ (.LO(la_data_out[95]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _111_ (.LO(la_data_out[96]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _112_ (.LO(la_data_out[97]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _113_ (.LO(la_data_out[98]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _114_ (.LO(la_data_out[99]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _115_ (.LO(la_data_out[100]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _116_ (.LO(la_data_out[101]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _117_ (.LO(la_data_out[102]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _118_ (.LO(la_data_out[103]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _119_ (.LO(la_data_out[104]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _120_ (.LO(la_data_out[105]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _121_ (.LO(la_data_out[106]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _122_ (.LO(la_data_out[107]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _123_ (.LO(la_data_out[108]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _124_ (.LO(la_data_out[109]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _125_ (.LO(la_data_out[110]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _126_ (.LO(la_data_out[111]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _127_ (.LO(la_data_out[112]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _128_ (.LO(la_data_out[113]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _129_ (.LO(la_data_out[114]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _130_ (.LO(la_data_out[115]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _131_ (.LO(la_data_out[116]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _132_ (.LO(la_data_out[117]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _133_ (.LO(la_data_out[118]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _134_ (.LO(la_data_out[119]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _135_ (.LO(la_data_out[120]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _136_ (.LO(la_data_out[121]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _137_ (.LO(la_data_out[122]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _138_ (.LO(la_data_out[123]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _139_ (.LO(la_data_out[124]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _140_ (.LO(la_data_out[125]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _141_ (.LO(la_data_out[126]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _142_ (.LO(la_data_out[127]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _143_ (.LO(io_out[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _144_ (.LO(io_out[37]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _145_ (.LO(io_oeb[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _146_ (.LO(io_oeb[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _147_ (.LO(io_oeb[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _148_ (.LO(io_oeb[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _149_ (.LO(io_oeb[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _150_ (.LO(io_oeb[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _151_ (.LO(io_oeb[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _152_ (.LO(io_oeb[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _153_ (.LO(io_oeb[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _154_ (.LO(io_oeb[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _155_ (.LO(io_oeb[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _156_ (.LO(io_oeb[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _157_ (.LO(io_oeb[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _158_ (.LO(io_oeb[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _159_ (.LO(io_oeb[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _160_ (.LO(io_oeb[16]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _161_ (.LO(io_oeb[17]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _162_ (.LO(io_oeb[18]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _163_ (.LO(io_oeb[19]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _164_ (.LO(io_oeb[20]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _165_ (.LO(io_oeb[21]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _166_ (.LO(io_oeb[22]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _167_ (.LO(io_oeb[23]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _168_ (.LO(io_oeb[24]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _169_ (.LO(io_oeb[25]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _170_ (.LO(io_oeb[26]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _171_ (.LO(io_oeb[27]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _172_ (.LO(io_oeb[28]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _173_ (.LO(io_oeb[29]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _174_ (.LO(io_oeb[30]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _175_ (.LO(io_oeb[31]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _176_ (.LO(_003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _177_ (.LO(_004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _178_ (.LO(_005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _179_ (.LO(_006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _180_ (.LO(_007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _181_ (.A(\u_core.sdr_den_n ),
    .X(io_oeb[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _182_ (.A(io_oeb[35]),
    .X(io_oeb[32]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _183_ (.A(io_oeb[35]),
    .X(io_oeb[33]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _184_ (.A(io_oeb[35]),
    .X(io_oeb[34]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_4 _185_ (.A(\u_core.sdr_dqm ),
    .X(io_out[23]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_4 _186_ (.A(\u_core.sdr_we_n ),
    .X(io_out[24]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_4 _187_ (.A(\u_core.sdr_cas_n ),
    .X(io_out[25]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_4 _188_ (.A(\u_core.sdr_ras_n ),
    .X(io_out[26]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _189_ (.A(\u_core.sdr_cs_n ),
    .X(io_out[27]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_4 _190_ (.A(\u_core.sdr_cke ),
    .X(io_out[28]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _191_ (.A(\u_core.sdram_clk ),
    .X(io_out[29]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _192_ (.A(\u_core.spim_clk ),
    .X(io_out[30]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _193_ (.A(\u_core.spim_csn ),
    .X(io_out[31]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _194_ (.A(\u_core.spim_sdo0 ),
    .X(io_out[32]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _195_ (.A(\u_core.spim_sdo1 ),
    .X(io_out[33]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _196_ (.A(\u_core.spim_sdo2 ),
    .X(io_out[34]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _197_ (.A(\u_core.spim_sdo3 ),
    .X(io_out[35]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 glbl_cfg \u_core.u_glbl_cfg  (.cfg_sdr_en(\u_core.cfg_sdr_en ),
    .cpu_rst_n(\u_core.cpu_rst_n ),
    .mclk(wb_clk_i),
    .reg_ack(\u_core.wbd_glbl_ack_i ),
    .reg_cs(\u_core.wbd_glbl_stb_o ),
    .reg_wr(\u_core.wbd_glbl_we_o ),
    .reset_n(\u_core.wb_rst_n ),
    .sdr_init_done(\u_core.sdr_init_done ),
    .sdram_clk(\u_core.sdram_clk ),
    .sdram_rst_n(\u_core.sdram_rst_n ),
    .soft_irq(\u_core.soft_irq ),
    .spi_rst_n(\u_core.spi_rst_n ),
    .VPWR(vccd1),
    .VGND(vssd1),
    .cfg_colbits({\u_core.cfg_colbits[1] ,
    \u_core.cfg_colbits[0] }),
    .cfg_req_depth({\u_core.cfg_req_depth[1] ,
    \u_core.cfg_req_depth[0] }),
    .cfg_sdr_cas({\u_core.cfg_sdr_cas[2] ,
    \u_core.cfg_sdr_cas[1] ,
    \u_core.cfg_sdr_cas[0] }),
    .cfg_sdr_mode_reg({\u_core.cfg_sdr_mode_reg[12] ,
    \u_core.cfg_sdr_mode_reg[11] ,
    \u_core.cfg_sdr_mode_reg[10] ,
    \u_core.cfg_sdr_mode_reg[9] ,
    \u_core.cfg_sdr_mode_reg[8] ,
    \u_core.cfg_sdr_mode_reg[7] ,
    \u_core.cfg_sdr_mode_reg[6] ,
    \u_core.cfg_sdr_mode_reg[5] ,
    \u_core.cfg_sdr_mode_reg[4] ,
    \u_core.cfg_sdr_mode_reg[3] ,
    \u_core.cfg_sdr_mode_reg[2] ,
    \u_core.cfg_sdr_mode_reg[1] ,
    \u_core.cfg_sdr_mode_reg[0] }),
    .cfg_sdr_rfmax({\u_core.cfg_sdr_rfmax[2] ,
    \u_core.cfg_sdr_rfmax[1] ,
    \u_core.cfg_sdr_rfmax[0] }),
    .cfg_sdr_rfsh({\u_core.cfg_sdr_rfsh[11] ,
    \u_core.cfg_sdr_rfsh[10] ,
    \u_core.cfg_sdr_rfsh[9] ,
    \u_core.cfg_sdr_rfsh[8] ,
    \u_core.cfg_sdr_rfsh[7] ,
    \u_core.cfg_sdr_rfsh[6] ,
    \u_core.cfg_sdr_rfsh[5] ,
    \u_core.cfg_sdr_rfsh[4] ,
    \u_core.cfg_sdr_rfsh[3] ,
    \u_core.cfg_sdr_rfsh[2] ,
    \u_core.cfg_sdr_rfsh[1] ,
    \u_core.cfg_sdr_rfsh[0] }),
    .cfg_sdr_tras_d({\u_core.cfg_sdr_tras_d[3] ,
    \u_core.cfg_sdr_tras_d[2] ,
    \u_core.cfg_sdr_tras_d[1] ,
    \u_core.cfg_sdr_tras_d[0] }),
    .cfg_sdr_trcar_d({\u_core.cfg_sdr_trcar_d[3] ,
    \u_core.cfg_sdr_trcar_d[2] ,
    \u_core.cfg_sdr_trcar_d[1] ,
    \u_core.cfg_sdr_trcar_d[0] }),
    .cfg_sdr_trcd_d({\u_core.cfg_sdr_trcd_d[3] ,
    \u_core.cfg_sdr_trcd_d[2] ,
    \u_core.cfg_sdr_trcd_d[1] ,
    \u_core.cfg_sdr_trcd_d[0] }),
    .cfg_sdr_trp_d({\u_core.cfg_sdr_trp_d[3] ,
    \u_core.cfg_sdr_trp_d[2] ,
    \u_core.cfg_sdr_trp_d[1] ,
    \u_core.cfg_sdr_trp_d[0] }),
    .cfg_sdr_twr_d({\u_core.cfg_sdr_twr_d[3] ,
    \u_core.cfg_sdr_twr_d[2] ,
    \u_core.cfg_sdr_twr_d[1] ,
    \u_core.cfg_sdr_twr_d[0] }),
    .cfg_sdr_width({\u_core.cfg_sdr_width[1] ,
    \u_core.cfg_sdr_width[0] }),
    .device_idcode({_NC1,
    _NC2,
    _NC3,
    _NC4,
    _NC5,
    _NC6,
    _NC7,
    _NC8,
    _NC9,
    _NC10,
    _NC11,
    _NC12,
    _NC13,
    _NC14,
    _NC15,
    _NC16,
    _NC17,
    _NC18,
    _NC19,
    _NC20,
    _NC21,
    _NC22,
    _NC23,
    _NC24,
    _NC25,
    _NC26,
    _NC27,
    _NC28,
    _NC29,
    _NC30,
    _NC31,
    _NC32}),
    .fuse_mhartid({\u_core.fuse_mhartid[31] ,
    \u_core.fuse_mhartid[30] ,
    \u_core.fuse_mhartid[29] ,
    \u_core.fuse_mhartid[28] ,
    \u_core.fuse_mhartid[27] ,
    \u_core.fuse_mhartid[26] ,
    \u_core.fuse_mhartid[25] ,
    \u_core.fuse_mhartid[24] ,
    \u_core.fuse_mhartid[23] ,
    \u_core.fuse_mhartid[22] ,
    \u_core.fuse_mhartid[21] ,
    \u_core.fuse_mhartid[20] ,
    \u_core.fuse_mhartid[19] ,
    \u_core.fuse_mhartid[18] ,
    \u_core.fuse_mhartid[17] ,
    \u_core.fuse_mhartid[16] ,
    \u_core.fuse_mhartid[15] ,
    \u_core.fuse_mhartid[14] ,
    \u_core.fuse_mhartid[13] ,
    \u_core.fuse_mhartid[12] ,
    \u_core.fuse_mhartid[11] ,
    \u_core.fuse_mhartid[10] ,
    \u_core.fuse_mhartid[9] ,
    \u_core.fuse_mhartid[8] ,
    \u_core.fuse_mhartid[7] ,
    \u_core.fuse_mhartid[6] ,
    \u_core.fuse_mhartid[5] ,
    \u_core.fuse_mhartid[4] ,
    \u_core.fuse_mhartid[3] ,
    \u_core.fuse_mhartid[2] ,
    \u_core.fuse_mhartid[1] ,
    \u_core.fuse_mhartid[0] }),
    .irq_lines({\u_core.irq_lines[15] ,
    \u_core.irq_lines[14] ,
    \u_core.irq_lines[13] ,
    \u_core.irq_lines[12] ,
    \u_core.irq_lines[11] ,
    \u_core.irq_lines[10] ,
    \u_core.irq_lines[9] ,
    \u_core.irq_lines[8] ,
    \u_core.irq_lines[7] ,
    \u_core.irq_lines[6] ,
    \u_core.irq_lines[5] ,
    \u_core.irq_lines[4] ,
    \u_core.irq_lines[3] ,
    \u_core.irq_lines[2] ,
    \u_core.irq_lines[1] ,
    \u_core.irq_lines[0] }),
    .reg_addr({\u_core.wbd_glbl_adr_o[5] ,
    \u_core.wbd_glbl_adr_o[4] ,
    \u_core.wbd_glbl_adr_o[3] ,
    \u_core.wbd_glbl_adr_o[2] }),
    .reg_be({\u_core.wbd_glbl_sel_o[3] ,
    \u_core.wbd_glbl_sel_o[2] ,
    \u_core.wbd_glbl_sel_o[1] ,
    \u_core.wbd_glbl_sel_o[0] }),
    .reg_rdata({\u_core.wbd_glbl_dat_i[31] ,
    \u_core.wbd_glbl_dat_i[30] ,
    \u_core.wbd_glbl_dat_i[29] ,
    \u_core.wbd_glbl_dat_i[28] ,
    \u_core.wbd_glbl_dat_i[27] ,
    \u_core.wbd_glbl_dat_i[26] ,
    \u_core.wbd_glbl_dat_i[25] ,
    \u_core.wbd_glbl_dat_i[24] ,
    \u_core.wbd_glbl_dat_i[23] ,
    \u_core.wbd_glbl_dat_i[22] ,
    \u_core.wbd_glbl_dat_i[21] ,
    \u_core.wbd_glbl_dat_i[20] ,
    \u_core.wbd_glbl_dat_i[19] ,
    \u_core.wbd_glbl_dat_i[18] ,
    \u_core.wbd_glbl_dat_i[17] ,
    \u_core.wbd_glbl_dat_i[16] ,
    \u_core.wbd_glbl_dat_i[15] ,
    \u_core.wbd_glbl_dat_i[14] ,
    \u_core.wbd_glbl_dat_i[13] ,
    \u_core.wbd_glbl_dat_i[12] ,
    \u_core.wbd_glbl_dat_i[11] ,
    \u_core.wbd_glbl_dat_i[10] ,
    \u_core.wbd_glbl_dat_i[9] ,
    \u_core.wbd_glbl_dat_i[8] ,
    \u_core.wbd_glbl_dat_i[7] ,
    \u_core.wbd_glbl_dat_i[6] ,
    \u_core.wbd_glbl_dat_i[5] ,
    \u_core.wbd_glbl_dat_i[4] ,
    \u_core.wbd_glbl_dat_i[3] ,
    \u_core.wbd_glbl_dat_i[2] ,
    \u_core.wbd_glbl_dat_i[1] ,
    \u_core.wbd_glbl_dat_i[0] }),
    .reg_wdata({\u_core.wbd_glbl_dat_o[31] ,
    \u_core.wbd_glbl_dat_o[30] ,
    \u_core.wbd_glbl_dat_o[29] ,
    \u_core.wbd_glbl_dat_o[28] ,
    \u_core.wbd_glbl_dat_o[27] ,
    \u_core.wbd_glbl_dat_o[26] ,
    \u_core.wbd_glbl_dat_o[25] ,
    \u_core.wbd_glbl_dat_o[24] ,
    \u_core.wbd_glbl_dat_o[23] ,
    \u_core.wbd_glbl_dat_o[22] ,
    \u_core.wbd_glbl_dat_o[21] ,
    \u_core.wbd_glbl_dat_o[20] ,
    \u_core.wbd_glbl_dat_o[19] ,
    \u_core.wbd_glbl_dat_o[18] ,
    \u_core.wbd_glbl_dat_o[17] ,
    \u_core.wbd_glbl_dat_o[16] ,
    \u_core.wbd_glbl_dat_o[15] ,
    \u_core.wbd_glbl_dat_o[14] ,
    \u_core.wbd_glbl_dat_o[13] ,
    \u_core.wbd_glbl_dat_o[12] ,
    \u_core.wbd_glbl_dat_o[11] ,
    \u_core.wbd_glbl_dat_o[10] ,
    \u_core.wbd_glbl_dat_o[9] ,
    \u_core.wbd_glbl_dat_o[8] ,
    \u_core.wbd_glbl_dat_o[7] ,
    \u_core.wbd_glbl_dat_o[6] ,
    \u_core.wbd_glbl_dat_o[5] ,
    \u_core.wbd_glbl_dat_o[4] ,
    \u_core.wbd_glbl_dat_o[3] ,
    \u_core.wbd_glbl_dat_o[2] ,
    \u_core.wbd_glbl_dat_o[1] ,
    \u_core.wbd_glbl_dat_o[0] }),
    .user_irq({user_irq[2],
    user_irq[1],
    user_irq[0]}));
 wb_interconnect \u_core.u_intercon  (.clk_i(wb_clk_i),
    .m0_wbd_ack_o(\u_core.wbd_riscv_imem_ack_o ),
    .m0_wbd_cyc_i(\u_core.wbd_riscv_imem_stb_i ),
    .m0_wbd_err_o(\u_core.wbd_riscv_imem_err_o ),
    .m0_wbd_stb_i(\u_core.wbd_riscv_imem_stb_i ),
    .m0_wbd_we_i(\u_core.wbd_riscv_imem_we_i ),
    .m1_wbd_ack_o(\u_core.wbd_riscv_dmem_ack_o ),
    .m1_wbd_cyc_i(\u_core.wbd_riscv_dmem_stb_i ),
    .m1_wbd_err_o(\u_core.wbd_riscv_dmem_err_o ),
    .m1_wbd_stb_i(\u_core.wbd_riscv_dmem_stb_i ),
    .m1_wbd_we_i(\u_core.wbd_riscv_dmem_we_i ),
    .m2_wbd_ack_o(wbs_ack_o),
    .m2_wbd_cyc_i(wbs_cyc_i),
    .m2_wbd_err_o(\u_core.wbd_ext_err_o ),
    .m2_wbd_stb_i(wbs_stb_i),
    .m2_wbd_we_i(wbs_we_i),
    .rst_n(\u_core.wb_rst_n ),
    .s0_wbd_ack_i(\u_core.wbd_spim_ack_i ),
    .s0_wbd_cyc_o(\u_core.wbd_spim_cyc_o ),
    .s0_wbd_err_i(_003_),
    .s0_wbd_stb_o(\u_core.wbd_spim_stb_o ),
    .s0_wbd_we_o(\u_core.wbd_spim_we_o ),
    .s1_wbd_ack_i(\u_core.wbd_sdram_ack_i ),
    .s1_wbd_cyc_o(\u_core.wbd_sdram_cyc_o ),
    .s1_wbd_err_i(_004_),
    .s1_wbd_stb_o(\u_core.wbd_sdram_stb_o ),
    .s1_wbd_we_o(\u_core.wbd_sdram_we_o ),
    .s2_wbd_ack_i(\u_core.wbd_glbl_ack_i ),
    .s2_wbd_cyc_o(\u_core.wbd_glbl_cyc_o ),
    .s2_wbd_err_i(_005_),
    .s2_wbd_stb_o(\u_core.wbd_glbl_stb_o ),
    .s2_wbd_we_o(\u_core.wbd_glbl_we_o ),
    .VPWR(vccd1),
    .VGND(vssd1),
    .m0_wbd_adr_i({\u_core.wbd_riscv_imem_adr_i[31] ,
    \u_core.wbd_riscv_imem_adr_i[30] ,
    \u_core.wbd_riscv_imem_adr_i[29] ,
    \u_core.wbd_riscv_imem_adr_i[28] ,
    \u_core.wbd_riscv_imem_adr_i[27] ,
    \u_core.wbd_riscv_imem_adr_i[26] ,
    \u_core.wbd_riscv_imem_adr_i[25] ,
    \u_core.wbd_riscv_imem_adr_i[24] ,
    \u_core.wbd_riscv_imem_adr_i[23] ,
    \u_core.wbd_riscv_imem_adr_i[22] ,
    \u_core.wbd_riscv_imem_adr_i[21] ,
    \u_core.wbd_riscv_imem_adr_i[20] ,
    \u_core.wbd_riscv_imem_adr_i[19] ,
    \u_core.wbd_riscv_imem_adr_i[18] ,
    \u_core.wbd_riscv_imem_adr_i[17] ,
    \u_core.wbd_riscv_imem_adr_i[16] ,
    \u_core.wbd_riscv_imem_adr_i[15] ,
    \u_core.wbd_riscv_imem_adr_i[14] ,
    \u_core.wbd_riscv_imem_adr_i[13] ,
    \u_core.wbd_riscv_imem_adr_i[12] ,
    \u_core.wbd_riscv_imem_adr_i[11] ,
    \u_core.wbd_riscv_imem_adr_i[10] ,
    \u_core.wbd_riscv_imem_adr_i[9] ,
    \u_core.wbd_riscv_imem_adr_i[8] ,
    \u_core.wbd_riscv_imem_adr_i[7] ,
    \u_core.wbd_riscv_imem_adr_i[6] ,
    \u_core.wbd_riscv_imem_adr_i[5] ,
    \u_core.wbd_riscv_imem_adr_i[4] ,
    \u_core.wbd_riscv_imem_adr_i[3] ,
    \u_core.wbd_riscv_imem_adr_i[2] ,
    \u_core.wbd_riscv_imem_adr_i[1] ,
    \u_core.wbd_riscv_imem_adr_i[0] }),
    .m0_wbd_dat_i({\u_core.wbd_riscv_imem_dat_i[31] ,
    \u_core.wbd_riscv_imem_dat_i[30] ,
    \u_core.wbd_riscv_imem_dat_i[29] ,
    \u_core.wbd_riscv_imem_dat_i[28] ,
    \u_core.wbd_riscv_imem_dat_i[27] ,
    \u_core.wbd_riscv_imem_dat_i[26] ,
    \u_core.wbd_riscv_imem_dat_i[25] ,
    \u_core.wbd_riscv_imem_dat_i[24] ,
    \u_core.wbd_riscv_imem_dat_i[23] ,
    \u_core.wbd_riscv_imem_dat_i[22] ,
    \u_core.wbd_riscv_imem_dat_i[21] ,
    \u_core.wbd_riscv_imem_dat_i[20] ,
    \u_core.wbd_riscv_imem_dat_i[19] ,
    \u_core.wbd_riscv_imem_dat_i[18] ,
    \u_core.wbd_riscv_imem_dat_i[17] ,
    \u_core.wbd_riscv_imem_dat_i[16] ,
    \u_core.wbd_riscv_imem_dat_i[15] ,
    \u_core.wbd_riscv_imem_dat_i[14] ,
    \u_core.wbd_riscv_imem_dat_i[13] ,
    \u_core.wbd_riscv_imem_dat_i[12] ,
    \u_core.wbd_riscv_imem_dat_i[11] ,
    \u_core.wbd_riscv_imem_dat_i[10] ,
    \u_core.wbd_riscv_imem_dat_i[9] ,
    \u_core.wbd_riscv_imem_dat_i[8] ,
    \u_core.wbd_riscv_imem_dat_i[7] ,
    \u_core.wbd_riscv_imem_dat_i[6] ,
    \u_core.wbd_riscv_imem_dat_i[5] ,
    \u_core.wbd_riscv_imem_dat_i[4] ,
    \u_core.wbd_riscv_imem_dat_i[3] ,
    \u_core.wbd_riscv_imem_dat_i[2] ,
    \u_core.wbd_riscv_imem_dat_i[1] ,
    \u_core.wbd_riscv_imem_dat_i[0] }),
    .m0_wbd_dat_o({\u_core.wbd_riscv_imem_dat_o[31] ,
    \u_core.wbd_riscv_imem_dat_o[30] ,
    \u_core.wbd_riscv_imem_dat_o[29] ,
    \u_core.wbd_riscv_imem_dat_o[28] ,
    \u_core.wbd_riscv_imem_dat_o[27] ,
    \u_core.wbd_riscv_imem_dat_o[26] ,
    \u_core.wbd_riscv_imem_dat_o[25] ,
    \u_core.wbd_riscv_imem_dat_o[24] ,
    \u_core.wbd_riscv_imem_dat_o[23] ,
    \u_core.wbd_riscv_imem_dat_o[22] ,
    \u_core.wbd_riscv_imem_dat_o[21] ,
    \u_core.wbd_riscv_imem_dat_o[20] ,
    \u_core.wbd_riscv_imem_dat_o[19] ,
    \u_core.wbd_riscv_imem_dat_o[18] ,
    \u_core.wbd_riscv_imem_dat_o[17] ,
    \u_core.wbd_riscv_imem_dat_o[16] ,
    \u_core.wbd_riscv_imem_dat_o[15] ,
    \u_core.wbd_riscv_imem_dat_o[14] ,
    \u_core.wbd_riscv_imem_dat_o[13] ,
    \u_core.wbd_riscv_imem_dat_o[12] ,
    \u_core.wbd_riscv_imem_dat_o[11] ,
    \u_core.wbd_riscv_imem_dat_o[10] ,
    \u_core.wbd_riscv_imem_dat_o[9] ,
    \u_core.wbd_riscv_imem_dat_o[8] ,
    \u_core.wbd_riscv_imem_dat_o[7] ,
    \u_core.wbd_riscv_imem_dat_o[6] ,
    \u_core.wbd_riscv_imem_dat_o[5] ,
    \u_core.wbd_riscv_imem_dat_o[4] ,
    \u_core.wbd_riscv_imem_dat_o[3] ,
    \u_core.wbd_riscv_imem_dat_o[2] ,
    \u_core.wbd_riscv_imem_dat_o[1] ,
    \u_core.wbd_riscv_imem_dat_o[0] }),
    .m0_wbd_sel_i({\u_core.wbd_riscv_imem_sel_i[3] ,
    \u_core.wbd_riscv_imem_sel_i[2] ,
    \u_core.wbd_riscv_imem_sel_i[1] ,
    \u_core.wbd_riscv_imem_sel_i[0] }),
    .m1_wbd_adr_i({\u_core.wbd_riscv_dmem_adr_i[31] ,
    \u_core.wbd_riscv_dmem_adr_i[30] ,
    \u_core.wbd_riscv_dmem_adr_i[29] ,
    \u_core.wbd_riscv_dmem_adr_i[28] ,
    \u_core.wbd_riscv_dmem_adr_i[27] ,
    \u_core.wbd_riscv_dmem_adr_i[26] ,
    \u_core.wbd_riscv_dmem_adr_i[25] ,
    \u_core.wbd_riscv_dmem_adr_i[24] ,
    \u_core.wbd_riscv_dmem_adr_i[23] ,
    \u_core.wbd_riscv_dmem_adr_i[22] ,
    \u_core.wbd_riscv_dmem_adr_i[21] ,
    \u_core.wbd_riscv_dmem_adr_i[20] ,
    \u_core.wbd_riscv_dmem_adr_i[19] ,
    \u_core.wbd_riscv_dmem_adr_i[18] ,
    \u_core.wbd_riscv_dmem_adr_i[17] ,
    \u_core.wbd_riscv_dmem_adr_i[16] ,
    \u_core.wbd_riscv_dmem_adr_i[15] ,
    \u_core.wbd_riscv_dmem_adr_i[14] ,
    \u_core.wbd_riscv_dmem_adr_i[13] ,
    \u_core.wbd_riscv_dmem_adr_i[12] ,
    \u_core.wbd_riscv_dmem_adr_i[11] ,
    \u_core.wbd_riscv_dmem_adr_i[10] ,
    \u_core.wbd_riscv_dmem_adr_i[9] ,
    \u_core.wbd_riscv_dmem_adr_i[8] ,
    \u_core.wbd_riscv_dmem_adr_i[7] ,
    \u_core.wbd_riscv_dmem_adr_i[6] ,
    \u_core.wbd_riscv_dmem_adr_i[5] ,
    \u_core.wbd_riscv_dmem_adr_i[4] ,
    \u_core.wbd_riscv_dmem_adr_i[3] ,
    \u_core.wbd_riscv_dmem_adr_i[2] ,
    \u_core.wbd_riscv_dmem_adr_i[1] ,
    \u_core.wbd_riscv_dmem_adr_i[0] }),
    .m1_wbd_dat_i({\u_core.wbd_riscv_dmem_dat_i[31] ,
    \u_core.wbd_riscv_dmem_dat_i[30] ,
    \u_core.wbd_riscv_dmem_dat_i[29] ,
    \u_core.wbd_riscv_dmem_dat_i[28] ,
    \u_core.wbd_riscv_dmem_dat_i[27] ,
    \u_core.wbd_riscv_dmem_dat_i[26] ,
    \u_core.wbd_riscv_dmem_dat_i[25] ,
    \u_core.wbd_riscv_dmem_dat_i[24] ,
    \u_core.wbd_riscv_dmem_dat_i[23] ,
    \u_core.wbd_riscv_dmem_dat_i[22] ,
    \u_core.wbd_riscv_dmem_dat_i[21] ,
    \u_core.wbd_riscv_dmem_dat_i[20] ,
    \u_core.wbd_riscv_dmem_dat_i[19] ,
    \u_core.wbd_riscv_dmem_dat_i[18] ,
    \u_core.wbd_riscv_dmem_dat_i[17] ,
    \u_core.wbd_riscv_dmem_dat_i[16] ,
    \u_core.wbd_riscv_dmem_dat_i[15] ,
    \u_core.wbd_riscv_dmem_dat_i[14] ,
    \u_core.wbd_riscv_dmem_dat_i[13] ,
    \u_core.wbd_riscv_dmem_dat_i[12] ,
    \u_core.wbd_riscv_dmem_dat_i[11] ,
    \u_core.wbd_riscv_dmem_dat_i[10] ,
    \u_core.wbd_riscv_dmem_dat_i[9] ,
    \u_core.wbd_riscv_dmem_dat_i[8] ,
    \u_core.wbd_riscv_dmem_dat_i[7] ,
    \u_core.wbd_riscv_dmem_dat_i[6] ,
    \u_core.wbd_riscv_dmem_dat_i[5] ,
    \u_core.wbd_riscv_dmem_dat_i[4] ,
    \u_core.wbd_riscv_dmem_dat_i[3] ,
    \u_core.wbd_riscv_dmem_dat_i[2] ,
    \u_core.wbd_riscv_dmem_dat_i[1] ,
    \u_core.wbd_riscv_dmem_dat_i[0] }),
    .m1_wbd_dat_o({\u_core.wbd_riscv_dmem_dat_o[31] ,
    \u_core.wbd_riscv_dmem_dat_o[30] ,
    \u_core.wbd_riscv_dmem_dat_o[29] ,
    \u_core.wbd_riscv_dmem_dat_o[28] ,
    \u_core.wbd_riscv_dmem_dat_o[27] ,
    \u_core.wbd_riscv_dmem_dat_o[26] ,
    \u_core.wbd_riscv_dmem_dat_o[25] ,
    \u_core.wbd_riscv_dmem_dat_o[24] ,
    \u_core.wbd_riscv_dmem_dat_o[23] ,
    \u_core.wbd_riscv_dmem_dat_o[22] ,
    \u_core.wbd_riscv_dmem_dat_o[21] ,
    \u_core.wbd_riscv_dmem_dat_o[20] ,
    \u_core.wbd_riscv_dmem_dat_o[19] ,
    \u_core.wbd_riscv_dmem_dat_o[18] ,
    \u_core.wbd_riscv_dmem_dat_o[17] ,
    \u_core.wbd_riscv_dmem_dat_o[16] ,
    \u_core.wbd_riscv_dmem_dat_o[15] ,
    \u_core.wbd_riscv_dmem_dat_o[14] ,
    \u_core.wbd_riscv_dmem_dat_o[13] ,
    \u_core.wbd_riscv_dmem_dat_o[12] ,
    \u_core.wbd_riscv_dmem_dat_o[11] ,
    \u_core.wbd_riscv_dmem_dat_o[10] ,
    \u_core.wbd_riscv_dmem_dat_o[9] ,
    \u_core.wbd_riscv_dmem_dat_o[8] ,
    \u_core.wbd_riscv_dmem_dat_o[7] ,
    \u_core.wbd_riscv_dmem_dat_o[6] ,
    \u_core.wbd_riscv_dmem_dat_o[5] ,
    \u_core.wbd_riscv_dmem_dat_o[4] ,
    \u_core.wbd_riscv_dmem_dat_o[3] ,
    \u_core.wbd_riscv_dmem_dat_o[2] ,
    \u_core.wbd_riscv_dmem_dat_o[1] ,
    \u_core.wbd_riscv_dmem_dat_o[0] }),
    .m1_wbd_sel_i({\u_core.wbd_riscv_dmem_sel_i[3] ,
    \u_core.wbd_riscv_dmem_sel_i[2] ,
    \u_core.wbd_riscv_dmem_sel_i[1] ,
    \u_core.wbd_riscv_dmem_sel_i[0] }),
    .m2_wbd_adr_i({wbs_adr_i[31],
    wbs_adr_i[30],
    wbs_adr_i[29],
    wbs_adr_i[28],
    wbs_adr_i[27],
    wbs_adr_i[26],
    wbs_adr_i[25],
    wbs_adr_i[24],
    wbs_adr_i[23],
    wbs_adr_i[22],
    wbs_adr_i[21],
    wbs_adr_i[20],
    wbs_adr_i[19],
    wbs_adr_i[18],
    wbs_adr_i[17],
    wbs_adr_i[16],
    wbs_adr_i[15],
    wbs_adr_i[14],
    wbs_adr_i[13],
    wbs_adr_i[12],
    wbs_adr_i[11],
    wbs_adr_i[10],
    wbs_adr_i[9],
    wbs_adr_i[8],
    wbs_adr_i[7],
    wbs_adr_i[6],
    wbs_adr_i[5],
    wbs_adr_i[4],
    wbs_adr_i[3],
    wbs_adr_i[2],
    wbs_adr_i[1],
    wbs_adr_i[0]}),
    .m2_wbd_dat_i({wbs_dat_i[31],
    wbs_dat_i[30],
    wbs_dat_i[29],
    wbs_dat_i[28],
    wbs_dat_i[27],
    wbs_dat_i[26],
    wbs_dat_i[25],
    wbs_dat_i[24],
    wbs_dat_i[23],
    wbs_dat_i[22],
    wbs_dat_i[21],
    wbs_dat_i[20],
    wbs_dat_i[19],
    wbs_dat_i[18],
    wbs_dat_i[17],
    wbs_dat_i[16],
    wbs_dat_i[15],
    wbs_dat_i[14],
    wbs_dat_i[13],
    wbs_dat_i[12],
    wbs_dat_i[11],
    wbs_dat_i[10],
    wbs_dat_i[9],
    wbs_dat_i[8],
    wbs_dat_i[7],
    wbs_dat_i[6],
    wbs_dat_i[5],
    wbs_dat_i[4],
    wbs_dat_i[3],
    wbs_dat_i[2],
    wbs_dat_i[1],
    wbs_dat_i[0]}),
    .m2_wbd_dat_o({wbs_dat_o[31],
    wbs_dat_o[30],
    wbs_dat_o[29],
    wbs_dat_o[28],
    wbs_dat_o[27],
    wbs_dat_o[26],
    wbs_dat_o[25],
    wbs_dat_o[24],
    wbs_dat_o[23],
    wbs_dat_o[22],
    wbs_dat_o[21],
    wbs_dat_o[20],
    wbs_dat_o[19],
    wbs_dat_o[18],
    wbs_dat_o[17],
    wbs_dat_o[16],
    wbs_dat_o[15],
    wbs_dat_o[14],
    wbs_dat_o[13],
    wbs_dat_o[12],
    wbs_dat_o[11],
    wbs_dat_o[10],
    wbs_dat_o[9],
    wbs_dat_o[8],
    wbs_dat_o[7],
    wbs_dat_o[6],
    wbs_dat_o[5],
    wbs_dat_o[4],
    wbs_dat_o[3],
    wbs_dat_o[2],
    wbs_dat_o[1],
    wbs_dat_o[0]}),
    .m2_wbd_sel_i({wbs_sel_i[3],
    wbs_sel_i[2],
    wbs_sel_i[1],
    wbs_sel_i[0]}),
    .s0_wbd_adr_o({\u_core.wbd_spim_adr_o[31] ,
    \u_core.wbd_spim_adr_o[30] ,
    \u_core.wbd_spim_adr_o[29] ,
    \u_core.wbd_spim_adr_o[28] ,
    \u_core.wbd_spim_adr_o[27] ,
    \u_core.wbd_spim_adr_o[26] ,
    \u_core.wbd_spim_adr_o[25] ,
    \u_core.wbd_spim_adr_o[24] ,
    \u_core.wbd_spim_adr_o[23] ,
    \u_core.wbd_spim_adr_o[22] ,
    \u_core.wbd_spim_adr_o[21] ,
    \u_core.wbd_spim_adr_o[20] ,
    \u_core.wbd_spim_adr_o[19] ,
    \u_core.wbd_spim_adr_o[18] ,
    \u_core.wbd_spim_adr_o[17] ,
    \u_core.wbd_spim_adr_o[16] ,
    \u_core.wbd_spim_adr_o[15] ,
    \u_core.wbd_spim_adr_o[14] ,
    \u_core.wbd_spim_adr_o[13] ,
    \u_core.wbd_spim_adr_o[12] ,
    \u_core.wbd_spim_adr_o[11] ,
    \u_core.wbd_spim_adr_o[10] ,
    \u_core.wbd_spim_adr_o[9] ,
    \u_core.wbd_spim_adr_o[8] ,
    \u_core.wbd_spim_adr_o[7] ,
    \u_core.wbd_spim_adr_o[6] ,
    \u_core.wbd_spim_adr_o[5] ,
    \u_core.wbd_spim_adr_o[4] ,
    \u_core.wbd_spim_adr_o[3] ,
    \u_core.wbd_spim_adr_o[2] ,
    \u_core.wbd_spim_adr_o[1] ,
    \u_core.wbd_spim_adr_o[0] }),
    .s0_wbd_dat_i({\u_core.wbd_spim_dat_i[31] ,
    \u_core.wbd_spim_dat_i[30] ,
    \u_core.wbd_spim_dat_i[29] ,
    \u_core.wbd_spim_dat_i[28] ,
    \u_core.wbd_spim_dat_i[27] ,
    \u_core.wbd_spim_dat_i[26] ,
    \u_core.wbd_spim_dat_i[25] ,
    \u_core.wbd_spim_dat_i[24] ,
    \u_core.wbd_spim_dat_i[23] ,
    \u_core.wbd_spim_dat_i[22] ,
    \u_core.wbd_spim_dat_i[21] ,
    \u_core.wbd_spim_dat_i[20] ,
    \u_core.wbd_spim_dat_i[19] ,
    \u_core.wbd_spim_dat_i[18] ,
    \u_core.wbd_spim_dat_i[17] ,
    \u_core.wbd_spim_dat_i[16] ,
    \u_core.wbd_spim_dat_i[15] ,
    \u_core.wbd_spim_dat_i[14] ,
    \u_core.wbd_spim_dat_i[13] ,
    \u_core.wbd_spim_dat_i[12] ,
    \u_core.wbd_spim_dat_i[11] ,
    \u_core.wbd_spim_dat_i[10] ,
    \u_core.wbd_spim_dat_i[9] ,
    \u_core.wbd_spim_dat_i[8] ,
    \u_core.wbd_spim_dat_i[7] ,
    \u_core.wbd_spim_dat_i[6] ,
    \u_core.wbd_spim_dat_i[5] ,
    \u_core.wbd_spim_dat_i[4] ,
    \u_core.wbd_spim_dat_i[3] ,
    \u_core.wbd_spim_dat_i[2] ,
    \u_core.wbd_spim_dat_i[1] ,
    \u_core.wbd_spim_dat_i[0] }),
    .s0_wbd_dat_o({\u_core.wbd_spim_dat_o[31] ,
    \u_core.wbd_spim_dat_o[30] ,
    \u_core.wbd_spim_dat_o[29] ,
    \u_core.wbd_spim_dat_o[28] ,
    \u_core.wbd_spim_dat_o[27] ,
    \u_core.wbd_spim_dat_o[26] ,
    \u_core.wbd_spim_dat_o[25] ,
    \u_core.wbd_spim_dat_o[24] ,
    \u_core.wbd_spim_dat_o[23] ,
    \u_core.wbd_spim_dat_o[22] ,
    \u_core.wbd_spim_dat_o[21] ,
    \u_core.wbd_spim_dat_o[20] ,
    \u_core.wbd_spim_dat_o[19] ,
    \u_core.wbd_spim_dat_o[18] ,
    \u_core.wbd_spim_dat_o[17] ,
    \u_core.wbd_spim_dat_o[16] ,
    \u_core.wbd_spim_dat_o[15] ,
    \u_core.wbd_spim_dat_o[14] ,
    \u_core.wbd_spim_dat_o[13] ,
    \u_core.wbd_spim_dat_o[12] ,
    \u_core.wbd_spim_dat_o[11] ,
    \u_core.wbd_spim_dat_o[10] ,
    \u_core.wbd_spim_dat_o[9] ,
    \u_core.wbd_spim_dat_o[8] ,
    \u_core.wbd_spim_dat_o[7] ,
    \u_core.wbd_spim_dat_o[6] ,
    \u_core.wbd_spim_dat_o[5] ,
    \u_core.wbd_spim_dat_o[4] ,
    \u_core.wbd_spim_dat_o[3] ,
    \u_core.wbd_spim_dat_o[2] ,
    \u_core.wbd_spim_dat_o[1] ,
    \u_core.wbd_spim_dat_o[0] }),
    .s0_wbd_sel_o({\u_core.wbd_spim_sel_o[3] ,
    \u_core.wbd_spim_sel_o[2] ,
    \u_core.wbd_spim_sel_o[1] ,
    \u_core.wbd_spim_sel_o[0] }),
    .s1_wbd_adr_o({\u_core.wbd_sdram_adr_o[31] ,
    \u_core.wbd_sdram_adr_o[30] ,
    \u_core.wbd_sdram_adr_o[29] ,
    \u_core.wbd_sdram_adr_o[28] ,
    \u_core.wbd_sdram_adr_o[27] ,
    \u_core.wbd_sdram_adr_o[26] ,
    \u_core.wbd_sdram_adr_o[25] ,
    \u_core.wbd_sdram_adr_o[24] ,
    \u_core.wbd_sdram_adr_o[23] ,
    \u_core.wbd_sdram_adr_o[22] ,
    \u_core.wbd_sdram_adr_o[21] ,
    \u_core.wbd_sdram_adr_o[20] ,
    \u_core.wbd_sdram_adr_o[19] ,
    \u_core.wbd_sdram_adr_o[18] ,
    \u_core.wbd_sdram_adr_o[17] ,
    \u_core.wbd_sdram_adr_o[16] ,
    \u_core.wbd_sdram_adr_o[15] ,
    \u_core.wbd_sdram_adr_o[14] ,
    \u_core.wbd_sdram_adr_o[13] ,
    \u_core.wbd_sdram_adr_o[12] ,
    \u_core.wbd_sdram_adr_o[11] ,
    \u_core.wbd_sdram_adr_o[10] ,
    \u_core.wbd_sdram_adr_o[9] ,
    \u_core.wbd_sdram_adr_o[8] ,
    \u_core.wbd_sdram_adr_o[7] ,
    \u_core.wbd_sdram_adr_o[6] ,
    \u_core.wbd_sdram_adr_o[5] ,
    \u_core.wbd_sdram_adr_o[4] ,
    \u_core.wbd_sdram_adr_o[3] ,
    \u_core.wbd_sdram_adr_o[2] ,
    \u_core.wbd_sdram_adr_o[1] ,
    \u_core.wbd_sdram_adr_o[0] }),
    .s1_wbd_dat_i({\u_core.wbd_sdram_dat_i[31] ,
    \u_core.wbd_sdram_dat_i[30] ,
    \u_core.wbd_sdram_dat_i[29] ,
    \u_core.wbd_sdram_dat_i[28] ,
    \u_core.wbd_sdram_dat_i[27] ,
    \u_core.wbd_sdram_dat_i[26] ,
    \u_core.wbd_sdram_dat_i[25] ,
    \u_core.wbd_sdram_dat_i[24] ,
    \u_core.wbd_sdram_dat_i[23] ,
    \u_core.wbd_sdram_dat_i[22] ,
    \u_core.wbd_sdram_dat_i[21] ,
    \u_core.wbd_sdram_dat_i[20] ,
    \u_core.wbd_sdram_dat_i[19] ,
    \u_core.wbd_sdram_dat_i[18] ,
    \u_core.wbd_sdram_dat_i[17] ,
    \u_core.wbd_sdram_dat_i[16] ,
    \u_core.wbd_sdram_dat_i[15] ,
    \u_core.wbd_sdram_dat_i[14] ,
    \u_core.wbd_sdram_dat_i[13] ,
    \u_core.wbd_sdram_dat_i[12] ,
    \u_core.wbd_sdram_dat_i[11] ,
    \u_core.wbd_sdram_dat_i[10] ,
    \u_core.wbd_sdram_dat_i[9] ,
    \u_core.wbd_sdram_dat_i[8] ,
    \u_core.wbd_sdram_dat_i[7] ,
    \u_core.wbd_sdram_dat_i[6] ,
    \u_core.wbd_sdram_dat_i[5] ,
    \u_core.wbd_sdram_dat_i[4] ,
    \u_core.wbd_sdram_dat_i[3] ,
    \u_core.wbd_sdram_dat_i[2] ,
    \u_core.wbd_sdram_dat_i[1] ,
    \u_core.wbd_sdram_dat_i[0] }),
    .s1_wbd_dat_o({\u_core.wbd_sdram_dat_o[31] ,
    \u_core.wbd_sdram_dat_o[30] ,
    \u_core.wbd_sdram_dat_o[29] ,
    \u_core.wbd_sdram_dat_o[28] ,
    \u_core.wbd_sdram_dat_o[27] ,
    \u_core.wbd_sdram_dat_o[26] ,
    \u_core.wbd_sdram_dat_o[25] ,
    \u_core.wbd_sdram_dat_o[24] ,
    \u_core.wbd_sdram_dat_o[23] ,
    \u_core.wbd_sdram_dat_o[22] ,
    \u_core.wbd_sdram_dat_o[21] ,
    \u_core.wbd_sdram_dat_o[20] ,
    \u_core.wbd_sdram_dat_o[19] ,
    \u_core.wbd_sdram_dat_o[18] ,
    \u_core.wbd_sdram_dat_o[17] ,
    \u_core.wbd_sdram_dat_o[16] ,
    \u_core.wbd_sdram_dat_o[15] ,
    \u_core.wbd_sdram_dat_o[14] ,
    \u_core.wbd_sdram_dat_o[13] ,
    \u_core.wbd_sdram_dat_o[12] ,
    \u_core.wbd_sdram_dat_o[11] ,
    \u_core.wbd_sdram_dat_o[10] ,
    \u_core.wbd_sdram_dat_o[9] ,
    \u_core.wbd_sdram_dat_o[8] ,
    \u_core.wbd_sdram_dat_o[7] ,
    \u_core.wbd_sdram_dat_o[6] ,
    \u_core.wbd_sdram_dat_o[5] ,
    \u_core.wbd_sdram_dat_o[4] ,
    \u_core.wbd_sdram_dat_o[3] ,
    \u_core.wbd_sdram_dat_o[2] ,
    \u_core.wbd_sdram_dat_o[1] ,
    \u_core.wbd_sdram_dat_o[0] }),
    .s1_wbd_sel_o({\u_core.wbd_sdram_sel_o[3] ,
    \u_core.wbd_sdram_sel_o[2] ,
    \u_core.wbd_sdram_sel_o[1] ,
    \u_core.wbd_sdram_sel_o[0] }),
    .s2_wbd_adr_o({\u_core.wbd_glbl_adr_o[31] ,
    \u_core.wbd_glbl_adr_o[30] ,
    \u_core.wbd_glbl_adr_o[29] ,
    \u_core.wbd_glbl_adr_o[28] ,
    \u_core.wbd_glbl_adr_o[27] ,
    \u_core.wbd_glbl_adr_o[26] ,
    \u_core.wbd_glbl_adr_o[25] ,
    \u_core.wbd_glbl_adr_o[24] ,
    \u_core.wbd_glbl_adr_o[23] ,
    \u_core.wbd_glbl_adr_o[22] ,
    \u_core.wbd_glbl_adr_o[21] ,
    \u_core.wbd_glbl_adr_o[20] ,
    \u_core.wbd_glbl_adr_o[19] ,
    \u_core.wbd_glbl_adr_o[18] ,
    \u_core.wbd_glbl_adr_o[17] ,
    \u_core.wbd_glbl_adr_o[16] ,
    \u_core.wbd_glbl_adr_o[15] ,
    \u_core.wbd_glbl_adr_o[14] ,
    \u_core.wbd_glbl_adr_o[13] ,
    \u_core.wbd_glbl_adr_o[12] ,
    \u_core.wbd_glbl_adr_o[11] ,
    \u_core.wbd_glbl_adr_o[10] ,
    \u_core.wbd_glbl_adr_o[9] ,
    \u_core.wbd_glbl_adr_o[8] ,
    \u_core.wbd_glbl_adr_o[7] ,
    \u_core.wbd_glbl_adr_o[6] ,
    \u_core.wbd_glbl_adr_o[5] ,
    \u_core.wbd_glbl_adr_o[4] ,
    \u_core.wbd_glbl_adr_o[3] ,
    \u_core.wbd_glbl_adr_o[2] ,
    \u_core.wbd_glbl_adr_o[1] ,
    \u_core.wbd_glbl_adr_o[0] }),
    .s2_wbd_dat_i({\u_core.wbd_glbl_dat_i[31] ,
    \u_core.wbd_glbl_dat_i[30] ,
    \u_core.wbd_glbl_dat_i[29] ,
    \u_core.wbd_glbl_dat_i[28] ,
    \u_core.wbd_glbl_dat_i[27] ,
    \u_core.wbd_glbl_dat_i[26] ,
    \u_core.wbd_glbl_dat_i[25] ,
    \u_core.wbd_glbl_dat_i[24] ,
    \u_core.wbd_glbl_dat_i[23] ,
    \u_core.wbd_glbl_dat_i[22] ,
    \u_core.wbd_glbl_dat_i[21] ,
    \u_core.wbd_glbl_dat_i[20] ,
    \u_core.wbd_glbl_dat_i[19] ,
    \u_core.wbd_glbl_dat_i[18] ,
    \u_core.wbd_glbl_dat_i[17] ,
    \u_core.wbd_glbl_dat_i[16] ,
    \u_core.wbd_glbl_dat_i[15] ,
    \u_core.wbd_glbl_dat_i[14] ,
    \u_core.wbd_glbl_dat_i[13] ,
    \u_core.wbd_glbl_dat_i[12] ,
    \u_core.wbd_glbl_dat_i[11] ,
    \u_core.wbd_glbl_dat_i[10] ,
    \u_core.wbd_glbl_dat_i[9] ,
    \u_core.wbd_glbl_dat_i[8] ,
    \u_core.wbd_glbl_dat_i[7] ,
    \u_core.wbd_glbl_dat_i[6] ,
    \u_core.wbd_glbl_dat_i[5] ,
    \u_core.wbd_glbl_dat_i[4] ,
    \u_core.wbd_glbl_dat_i[3] ,
    \u_core.wbd_glbl_dat_i[2] ,
    \u_core.wbd_glbl_dat_i[1] ,
    \u_core.wbd_glbl_dat_i[0] }),
    .s2_wbd_dat_o({\u_core.wbd_glbl_dat_o[31] ,
    \u_core.wbd_glbl_dat_o[30] ,
    \u_core.wbd_glbl_dat_o[29] ,
    \u_core.wbd_glbl_dat_o[28] ,
    \u_core.wbd_glbl_dat_o[27] ,
    \u_core.wbd_glbl_dat_o[26] ,
    \u_core.wbd_glbl_dat_o[25] ,
    \u_core.wbd_glbl_dat_o[24] ,
    \u_core.wbd_glbl_dat_o[23] ,
    \u_core.wbd_glbl_dat_o[22] ,
    \u_core.wbd_glbl_dat_o[21] ,
    \u_core.wbd_glbl_dat_o[20] ,
    \u_core.wbd_glbl_dat_o[19] ,
    \u_core.wbd_glbl_dat_o[18] ,
    \u_core.wbd_glbl_dat_o[17] ,
    \u_core.wbd_glbl_dat_o[16] ,
    \u_core.wbd_glbl_dat_o[15] ,
    \u_core.wbd_glbl_dat_o[14] ,
    \u_core.wbd_glbl_dat_o[13] ,
    \u_core.wbd_glbl_dat_o[12] ,
    \u_core.wbd_glbl_dat_o[11] ,
    \u_core.wbd_glbl_dat_o[10] ,
    \u_core.wbd_glbl_dat_o[9] ,
    \u_core.wbd_glbl_dat_o[8] ,
    \u_core.wbd_glbl_dat_o[7] ,
    \u_core.wbd_glbl_dat_o[6] ,
    \u_core.wbd_glbl_dat_o[5] ,
    \u_core.wbd_glbl_dat_o[4] ,
    \u_core.wbd_glbl_dat_o[3] ,
    \u_core.wbd_glbl_dat_o[2] ,
    \u_core.wbd_glbl_dat_o[1] ,
    \u_core.wbd_glbl_dat_o[0] }),
    .s2_wbd_sel_o({\u_core.wbd_glbl_sel_o[3] ,
    \u_core.wbd_glbl_sel_o[2] ,
    \u_core.wbd_glbl_sel_o[1] ,
    \u_core.wbd_glbl_sel_o[0] }));
 scr1_top_wb \u_core.u_riscv_top  (.clk(wb_clk_i),
    .cpu_rst_n(\u_core.cpu_rst_n ),
    .pwrup_rst_n(\u_core.wb_rst_n ),
    .rst_n(\u_core.wb_rst_n ),
    .rtc_clk(user_clock2),
    .soft_irq(\u_core.soft_irq ),
    .test_mode(_006_),
    .test_rst_n(_000_),
    .wbd_dmem_ack_i(\u_core.wbd_riscv_dmem_ack_o ),
    .wbd_dmem_err_i(\u_core.wbd_riscv_dmem_err_o ),
    .wbd_dmem_stb_o(\u_core.wbd_riscv_dmem_stb_i ),
    .wbd_dmem_we_o(\u_core.wbd_riscv_dmem_we_i ),
    .wbd_imem_ack_i(\u_core.wbd_riscv_imem_ack_o ),
    .wbd_imem_err_i(\u_core.wbd_riscv_imem_err_o ),
    .wbd_imem_stb_o(\u_core.wbd_riscv_imem_stb_i ),
    .wbd_imem_we_o(\u_core.wbd_riscv_imem_we_i ),
    .VPWR(vccd1),
    .VGND(vssd1),
    .fuse_mhartid({\u_core.fuse_mhartid[31] ,
    \u_core.fuse_mhartid[30] ,
    \u_core.fuse_mhartid[29] ,
    \u_core.fuse_mhartid[28] ,
    \u_core.fuse_mhartid[27] ,
    \u_core.fuse_mhartid[26] ,
    \u_core.fuse_mhartid[25] ,
    \u_core.fuse_mhartid[24] ,
    \u_core.fuse_mhartid[23] ,
    \u_core.fuse_mhartid[22] ,
    \u_core.fuse_mhartid[21] ,
    \u_core.fuse_mhartid[20] ,
    \u_core.fuse_mhartid[19] ,
    \u_core.fuse_mhartid[18] ,
    \u_core.fuse_mhartid[17] ,
    \u_core.fuse_mhartid[16] ,
    \u_core.fuse_mhartid[15] ,
    \u_core.fuse_mhartid[14] ,
    \u_core.fuse_mhartid[13] ,
    \u_core.fuse_mhartid[12] ,
    \u_core.fuse_mhartid[11] ,
    \u_core.fuse_mhartid[10] ,
    \u_core.fuse_mhartid[9] ,
    \u_core.fuse_mhartid[8] ,
    \u_core.fuse_mhartid[7] ,
    \u_core.fuse_mhartid[6] ,
    \u_core.fuse_mhartid[5] ,
    \u_core.fuse_mhartid[4] ,
    \u_core.fuse_mhartid[3] ,
    \u_core.fuse_mhartid[2] ,
    \u_core.fuse_mhartid[1] ,
    \u_core.fuse_mhartid[0] }),
    .irq_lines({\u_core.irq_lines[15] ,
    \u_core.irq_lines[14] ,
    \u_core.irq_lines[13] ,
    \u_core.irq_lines[12] ,
    \u_core.irq_lines[11] ,
    \u_core.irq_lines[10] ,
    \u_core.irq_lines[9] ,
    \u_core.irq_lines[8] ,
    \u_core.irq_lines[7] ,
    \u_core.irq_lines[6] ,
    \u_core.irq_lines[5] ,
    \u_core.irq_lines[4] ,
    \u_core.irq_lines[3] ,
    \u_core.irq_lines[2] ,
    \u_core.irq_lines[1] ,
    \u_core.irq_lines[0] }),
    .wbd_dmem_adr_o({\u_core.wbd_riscv_dmem_adr_i[31] ,
    \u_core.wbd_riscv_dmem_adr_i[30] ,
    \u_core.wbd_riscv_dmem_adr_i[29] ,
    \u_core.wbd_riscv_dmem_adr_i[28] ,
    \u_core.wbd_riscv_dmem_adr_i[27] ,
    \u_core.wbd_riscv_dmem_adr_i[26] ,
    \u_core.wbd_riscv_dmem_adr_i[25] ,
    \u_core.wbd_riscv_dmem_adr_i[24] ,
    \u_core.wbd_riscv_dmem_adr_i[23] ,
    \u_core.wbd_riscv_dmem_adr_i[22] ,
    \u_core.wbd_riscv_dmem_adr_i[21] ,
    \u_core.wbd_riscv_dmem_adr_i[20] ,
    \u_core.wbd_riscv_dmem_adr_i[19] ,
    \u_core.wbd_riscv_dmem_adr_i[18] ,
    \u_core.wbd_riscv_dmem_adr_i[17] ,
    \u_core.wbd_riscv_dmem_adr_i[16] ,
    \u_core.wbd_riscv_dmem_adr_i[15] ,
    \u_core.wbd_riscv_dmem_adr_i[14] ,
    \u_core.wbd_riscv_dmem_adr_i[13] ,
    \u_core.wbd_riscv_dmem_adr_i[12] ,
    \u_core.wbd_riscv_dmem_adr_i[11] ,
    \u_core.wbd_riscv_dmem_adr_i[10] ,
    \u_core.wbd_riscv_dmem_adr_i[9] ,
    \u_core.wbd_riscv_dmem_adr_i[8] ,
    \u_core.wbd_riscv_dmem_adr_i[7] ,
    \u_core.wbd_riscv_dmem_adr_i[6] ,
    \u_core.wbd_riscv_dmem_adr_i[5] ,
    \u_core.wbd_riscv_dmem_adr_i[4] ,
    \u_core.wbd_riscv_dmem_adr_i[3] ,
    \u_core.wbd_riscv_dmem_adr_i[2] ,
    \u_core.wbd_riscv_dmem_adr_i[1] ,
    \u_core.wbd_riscv_dmem_adr_i[0] }),
    .wbd_dmem_dat_i({\u_core.wbd_riscv_dmem_dat_o[31] ,
    \u_core.wbd_riscv_dmem_dat_o[30] ,
    \u_core.wbd_riscv_dmem_dat_o[29] ,
    \u_core.wbd_riscv_dmem_dat_o[28] ,
    \u_core.wbd_riscv_dmem_dat_o[27] ,
    \u_core.wbd_riscv_dmem_dat_o[26] ,
    \u_core.wbd_riscv_dmem_dat_o[25] ,
    \u_core.wbd_riscv_dmem_dat_o[24] ,
    \u_core.wbd_riscv_dmem_dat_o[23] ,
    \u_core.wbd_riscv_dmem_dat_o[22] ,
    \u_core.wbd_riscv_dmem_dat_o[21] ,
    \u_core.wbd_riscv_dmem_dat_o[20] ,
    \u_core.wbd_riscv_dmem_dat_o[19] ,
    \u_core.wbd_riscv_dmem_dat_o[18] ,
    \u_core.wbd_riscv_dmem_dat_o[17] ,
    \u_core.wbd_riscv_dmem_dat_o[16] ,
    \u_core.wbd_riscv_dmem_dat_o[15] ,
    \u_core.wbd_riscv_dmem_dat_o[14] ,
    \u_core.wbd_riscv_dmem_dat_o[13] ,
    \u_core.wbd_riscv_dmem_dat_o[12] ,
    \u_core.wbd_riscv_dmem_dat_o[11] ,
    \u_core.wbd_riscv_dmem_dat_o[10] ,
    \u_core.wbd_riscv_dmem_dat_o[9] ,
    \u_core.wbd_riscv_dmem_dat_o[8] ,
    \u_core.wbd_riscv_dmem_dat_o[7] ,
    \u_core.wbd_riscv_dmem_dat_o[6] ,
    \u_core.wbd_riscv_dmem_dat_o[5] ,
    \u_core.wbd_riscv_dmem_dat_o[4] ,
    \u_core.wbd_riscv_dmem_dat_o[3] ,
    \u_core.wbd_riscv_dmem_dat_o[2] ,
    \u_core.wbd_riscv_dmem_dat_o[1] ,
    \u_core.wbd_riscv_dmem_dat_o[0] }),
    .wbd_dmem_dat_o({\u_core.wbd_riscv_dmem_dat_i[31] ,
    \u_core.wbd_riscv_dmem_dat_i[30] ,
    \u_core.wbd_riscv_dmem_dat_i[29] ,
    \u_core.wbd_riscv_dmem_dat_i[28] ,
    \u_core.wbd_riscv_dmem_dat_i[27] ,
    \u_core.wbd_riscv_dmem_dat_i[26] ,
    \u_core.wbd_riscv_dmem_dat_i[25] ,
    \u_core.wbd_riscv_dmem_dat_i[24] ,
    \u_core.wbd_riscv_dmem_dat_i[23] ,
    \u_core.wbd_riscv_dmem_dat_i[22] ,
    \u_core.wbd_riscv_dmem_dat_i[21] ,
    \u_core.wbd_riscv_dmem_dat_i[20] ,
    \u_core.wbd_riscv_dmem_dat_i[19] ,
    \u_core.wbd_riscv_dmem_dat_i[18] ,
    \u_core.wbd_riscv_dmem_dat_i[17] ,
    \u_core.wbd_riscv_dmem_dat_i[16] ,
    \u_core.wbd_riscv_dmem_dat_i[15] ,
    \u_core.wbd_riscv_dmem_dat_i[14] ,
    \u_core.wbd_riscv_dmem_dat_i[13] ,
    \u_core.wbd_riscv_dmem_dat_i[12] ,
    \u_core.wbd_riscv_dmem_dat_i[11] ,
    \u_core.wbd_riscv_dmem_dat_i[10] ,
    \u_core.wbd_riscv_dmem_dat_i[9] ,
    \u_core.wbd_riscv_dmem_dat_i[8] ,
    \u_core.wbd_riscv_dmem_dat_i[7] ,
    \u_core.wbd_riscv_dmem_dat_i[6] ,
    \u_core.wbd_riscv_dmem_dat_i[5] ,
    \u_core.wbd_riscv_dmem_dat_i[4] ,
    \u_core.wbd_riscv_dmem_dat_i[3] ,
    \u_core.wbd_riscv_dmem_dat_i[2] ,
    \u_core.wbd_riscv_dmem_dat_i[1] ,
    \u_core.wbd_riscv_dmem_dat_i[0] }),
    .wbd_dmem_sel_o({\u_core.wbd_riscv_dmem_sel_i[3] ,
    \u_core.wbd_riscv_dmem_sel_i[2] ,
    \u_core.wbd_riscv_dmem_sel_i[1] ,
    \u_core.wbd_riscv_dmem_sel_i[0] }),
    .wbd_imem_adr_o({\u_core.wbd_riscv_imem_adr_i[31] ,
    \u_core.wbd_riscv_imem_adr_i[30] ,
    \u_core.wbd_riscv_imem_adr_i[29] ,
    \u_core.wbd_riscv_imem_adr_i[28] ,
    \u_core.wbd_riscv_imem_adr_i[27] ,
    \u_core.wbd_riscv_imem_adr_i[26] ,
    \u_core.wbd_riscv_imem_adr_i[25] ,
    \u_core.wbd_riscv_imem_adr_i[24] ,
    \u_core.wbd_riscv_imem_adr_i[23] ,
    \u_core.wbd_riscv_imem_adr_i[22] ,
    \u_core.wbd_riscv_imem_adr_i[21] ,
    \u_core.wbd_riscv_imem_adr_i[20] ,
    \u_core.wbd_riscv_imem_adr_i[19] ,
    \u_core.wbd_riscv_imem_adr_i[18] ,
    \u_core.wbd_riscv_imem_adr_i[17] ,
    \u_core.wbd_riscv_imem_adr_i[16] ,
    \u_core.wbd_riscv_imem_adr_i[15] ,
    \u_core.wbd_riscv_imem_adr_i[14] ,
    \u_core.wbd_riscv_imem_adr_i[13] ,
    \u_core.wbd_riscv_imem_adr_i[12] ,
    \u_core.wbd_riscv_imem_adr_i[11] ,
    \u_core.wbd_riscv_imem_adr_i[10] ,
    \u_core.wbd_riscv_imem_adr_i[9] ,
    \u_core.wbd_riscv_imem_adr_i[8] ,
    \u_core.wbd_riscv_imem_adr_i[7] ,
    \u_core.wbd_riscv_imem_adr_i[6] ,
    \u_core.wbd_riscv_imem_adr_i[5] ,
    \u_core.wbd_riscv_imem_adr_i[4] ,
    \u_core.wbd_riscv_imem_adr_i[3] ,
    \u_core.wbd_riscv_imem_adr_i[2] ,
    \u_core.wbd_riscv_imem_adr_i[1] ,
    \u_core.wbd_riscv_imem_adr_i[0] }),
    .wbd_imem_dat_i({\u_core.wbd_riscv_imem_dat_o[31] ,
    \u_core.wbd_riscv_imem_dat_o[30] ,
    \u_core.wbd_riscv_imem_dat_o[29] ,
    \u_core.wbd_riscv_imem_dat_o[28] ,
    \u_core.wbd_riscv_imem_dat_o[27] ,
    \u_core.wbd_riscv_imem_dat_o[26] ,
    \u_core.wbd_riscv_imem_dat_o[25] ,
    \u_core.wbd_riscv_imem_dat_o[24] ,
    \u_core.wbd_riscv_imem_dat_o[23] ,
    \u_core.wbd_riscv_imem_dat_o[22] ,
    \u_core.wbd_riscv_imem_dat_o[21] ,
    \u_core.wbd_riscv_imem_dat_o[20] ,
    \u_core.wbd_riscv_imem_dat_o[19] ,
    \u_core.wbd_riscv_imem_dat_o[18] ,
    \u_core.wbd_riscv_imem_dat_o[17] ,
    \u_core.wbd_riscv_imem_dat_o[16] ,
    \u_core.wbd_riscv_imem_dat_o[15] ,
    \u_core.wbd_riscv_imem_dat_o[14] ,
    \u_core.wbd_riscv_imem_dat_o[13] ,
    \u_core.wbd_riscv_imem_dat_o[12] ,
    \u_core.wbd_riscv_imem_dat_o[11] ,
    \u_core.wbd_riscv_imem_dat_o[10] ,
    \u_core.wbd_riscv_imem_dat_o[9] ,
    \u_core.wbd_riscv_imem_dat_o[8] ,
    \u_core.wbd_riscv_imem_dat_o[7] ,
    \u_core.wbd_riscv_imem_dat_o[6] ,
    \u_core.wbd_riscv_imem_dat_o[5] ,
    \u_core.wbd_riscv_imem_dat_o[4] ,
    \u_core.wbd_riscv_imem_dat_o[3] ,
    \u_core.wbd_riscv_imem_dat_o[2] ,
    \u_core.wbd_riscv_imem_dat_o[1] ,
    \u_core.wbd_riscv_imem_dat_o[0] }),
    .wbd_imem_dat_o({\u_core.wbd_riscv_imem_dat_i[31] ,
    \u_core.wbd_riscv_imem_dat_i[30] ,
    \u_core.wbd_riscv_imem_dat_i[29] ,
    \u_core.wbd_riscv_imem_dat_i[28] ,
    \u_core.wbd_riscv_imem_dat_i[27] ,
    \u_core.wbd_riscv_imem_dat_i[26] ,
    \u_core.wbd_riscv_imem_dat_i[25] ,
    \u_core.wbd_riscv_imem_dat_i[24] ,
    \u_core.wbd_riscv_imem_dat_i[23] ,
    \u_core.wbd_riscv_imem_dat_i[22] ,
    \u_core.wbd_riscv_imem_dat_i[21] ,
    \u_core.wbd_riscv_imem_dat_i[20] ,
    \u_core.wbd_riscv_imem_dat_i[19] ,
    \u_core.wbd_riscv_imem_dat_i[18] ,
    \u_core.wbd_riscv_imem_dat_i[17] ,
    \u_core.wbd_riscv_imem_dat_i[16] ,
    \u_core.wbd_riscv_imem_dat_i[15] ,
    \u_core.wbd_riscv_imem_dat_i[14] ,
    \u_core.wbd_riscv_imem_dat_i[13] ,
    \u_core.wbd_riscv_imem_dat_i[12] ,
    \u_core.wbd_riscv_imem_dat_i[11] ,
    \u_core.wbd_riscv_imem_dat_i[10] ,
    \u_core.wbd_riscv_imem_dat_i[9] ,
    \u_core.wbd_riscv_imem_dat_i[8] ,
    \u_core.wbd_riscv_imem_dat_i[7] ,
    \u_core.wbd_riscv_imem_dat_i[6] ,
    \u_core.wbd_riscv_imem_dat_i[5] ,
    \u_core.wbd_riscv_imem_dat_i[4] ,
    \u_core.wbd_riscv_imem_dat_i[3] ,
    \u_core.wbd_riscv_imem_dat_i[2] ,
    \u_core.wbd_riscv_imem_dat_i[1] ,
    \u_core.wbd_riscv_imem_dat_i[0] }),
    .wbd_imem_sel_o({\u_core.wbd_riscv_imem_sel_i[3] ,
    \u_core.wbd_riscv_imem_sel_i[2] ,
    \u_core.wbd_riscv_imem_sel_i[1] ,
    \u_core.wbd_riscv_imem_sel_i[0] }));
 sdrc_top \u_core.u_sdram_ctrl  (.cfg_sdr_en(\u_core.cfg_sdr_en ),
    .sdr_cas_n(\u_core.sdr_cas_n ),
    .sdr_cke(\u_core.sdr_cke ),
    .sdr_cs_n(\u_core.sdr_cs_n ),
    .sdr_den_n(\u_core.sdr_den_n ),
    .sdr_dqm(\u_core.sdr_dqm ),
    .sdr_init_done(\u_core.sdr_init_done ),
    .sdr_ras_n(\u_core.sdr_ras_n ),
    .sdr_we_n(\u_core.sdr_we_n ),
    .sdram_clk(\u_core.sdram_clk ),
    .sdram_pad_clk(io_in[29]),
    .sdram_resetn(\u_core.sdram_rst_n ),
    .wb_ack_o(\u_core.wbd_sdram_ack_i ),
    .wb_clk_i(wb_clk_i),
    .wb_cyc_i(\u_core.wbd_sdram_cyc_o ),
    .wb_rst_i(wb_rst_i),
    .wb_stb_i(\u_core.wbd_sdram_stb_o ),
    .wb_we_i(\u_core.wbd_sdram_we_o ),
    .VPWR(vccd1),
    .VGND(vssd1),
    .cfg_colbits({\u_core.cfg_colbits[1] ,
    \u_core.cfg_colbits[0] }),
    .cfg_req_depth({\u_core.cfg_req_depth[1] ,
    \u_core.cfg_req_depth[0] }),
    .cfg_sdr_cas({\u_core.cfg_sdr_cas[2] ,
    \u_core.cfg_sdr_cas[1] ,
    \u_core.cfg_sdr_cas[0] }),
    .cfg_sdr_mode_reg({\u_core.cfg_sdr_mode_reg[12] ,
    \u_core.cfg_sdr_mode_reg[11] ,
    \u_core.cfg_sdr_mode_reg[10] ,
    \u_core.cfg_sdr_mode_reg[9] ,
    \u_core.cfg_sdr_mode_reg[8] ,
    \u_core.cfg_sdr_mode_reg[7] ,
    \u_core.cfg_sdr_mode_reg[6] ,
    \u_core.cfg_sdr_mode_reg[5] ,
    \u_core.cfg_sdr_mode_reg[4] ,
    \u_core.cfg_sdr_mode_reg[3] ,
    \u_core.cfg_sdr_mode_reg[2] ,
    \u_core.cfg_sdr_mode_reg[1] ,
    \u_core.cfg_sdr_mode_reg[0] }),
    .cfg_sdr_rfmax({\u_core.cfg_sdr_rfmax[2] ,
    \u_core.cfg_sdr_rfmax[1] ,
    \u_core.cfg_sdr_rfmax[0] }),
    .cfg_sdr_rfsh({\u_core.cfg_sdr_rfsh[11] ,
    \u_core.cfg_sdr_rfsh[10] ,
    \u_core.cfg_sdr_rfsh[9] ,
    \u_core.cfg_sdr_rfsh[8] ,
    \u_core.cfg_sdr_rfsh[7] ,
    \u_core.cfg_sdr_rfsh[6] ,
    \u_core.cfg_sdr_rfsh[5] ,
    \u_core.cfg_sdr_rfsh[4] ,
    \u_core.cfg_sdr_rfsh[3] ,
    \u_core.cfg_sdr_rfsh[2] ,
    \u_core.cfg_sdr_rfsh[1] ,
    \u_core.cfg_sdr_rfsh[0] }),
    .cfg_sdr_tras_d({\u_core.cfg_sdr_tras_d[3] ,
    \u_core.cfg_sdr_tras_d[2] ,
    \u_core.cfg_sdr_tras_d[1] ,
    \u_core.cfg_sdr_tras_d[0] }),
    .cfg_sdr_trcar_d({\u_core.cfg_sdr_trcar_d[3] ,
    \u_core.cfg_sdr_trcar_d[2] ,
    \u_core.cfg_sdr_trcar_d[1] ,
    \u_core.cfg_sdr_trcar_d[0] }),
    .cfg_sdr_trcd_d({\u_core.cfg_sdr_trcd_d[3] ,
    \u_core.cfg_sdr_trcd_d[2] ,
    \u_core.cfg_sdr_trcd_d[1] ,
    \u_core.cfg_sdr_trcd_d[0] }),
    .cfg_sdr_trp_d({\u_core.cfg_sdr_trp_d[3] ,
    \u_core.cfg_sdr_trp_d[2] ,
    \u_core.cfg_sdr_trp_d[1] ,
    \u_core.cfg_sdr_trp_d[0] }),
    .cfg_sdr_twr_d({\u_core.cfg_sdr_twr_d[3] ,
    \u_core.cfg_sdr_twr_d[2] ,
    \u_core.cfg_sdr_twr_d[1] ,
    \u_core.cfg_sdr_twr_d[0] }),
    .cfg_sdr_width({\u_core.cfg_sdr_width[1] ,
    \u_core.cfg_sdr_width[0] }),
    .pad_sdr_din({io_in[7],
    io_in[6],
    io_in[5],
    io_in[4],
    io_in[3],
    io_in[2],
    io_in[1],
    io_in[0]}),
    .sdr_addr({io_out[20],
    io_out[19],
    io_out[18],
    io_out[17],
    io_out[16],
    io_out[15],
    io_out[14],
    io_out[13],
    io_out[12],
    io_out[11],
    io_out[10],
    io_out[9],
    io_out[8]}),
    .sdr_ba({io_out[22],
    io_out[21]}),
    .sdr_dout({io_out[7],
    io_out[6],
    io_out[5],
    io_out[4],
    io_out[3],
    io_out[2],
    io_out[1],
    io_out[0]}),
    .wb_addr_i({\u_core.wbd_sdram_adr_o[31] ,
    \u_core.wbd_sdram_adr_o[30] ,
    \u_core.wbd_sdram_adr_o[29] ,
    \u_core.wbd_sdram_adr_o[28] ,
    \u_core.wbd_sdram_adr_o[27] ,
    \u_core.wbd_sdram_adr_o[26] ,
    \u_core.wbd_sdram_adr_o[25] ,
    \u_core.wbd_sdram_adr_o[24] ,
    \u_core.wbd_sdram_adr_o[23] ,
    \u_core.wbd_sdram_adr_o[22] ,
    \u_core.wbd_sdram_adr_o[21] ,
    \u_core.wbd_sdram_adr_o[20] ,
    \u_core.wbd_sdram_adr_o[19] ,
    \u_core.wbd_sdram_adr_o[18] ,
    \u_core.wbd_sdram_adr_o[17] ,
    \u_core.wbd_sdram_adr_o[16] ,
    \u_core.wbd_sdram_adr_o[15] ,
    \u_core.wbd_sdram_adr_o[14] ,
    \u_core.wbd_sdram_adr_o[13] ,
    \u_core.wbd_sdram_adr_o[12] ,
    \u_core.wbd_sdram_adr_o[11] ,
    \u_core.wbd_sdram_adr_o[10] ,
    \u_core.wbd_sdram_adr_o[9] ,
    \u_core.wbd_sdram_adr_o[8] ,
    \u_core.wbd_sdram_adr_o[7] ,
    \u_core.wbd_sdram_adr_o[6] ,
    \u_core.wbd_sdram_adr_o[5] ,
    \u_core.wbd_sdram_adr_o[4] ,
    \u_core.wbd_sdram_adr_o[3] ,
    \u_core.wbd_sdram_adr_o[2] ,
    \u_core.wbd_sdram_adr_o[1] ,
    \u_core.wbd_sdram_adr_o[0] }),
    .wb_cti_i({_002_,
    _001_,
    _007_}),
    .wb_dat_i({\u_core.wbd_sdram_dat_o[31] ,
    \u_core.wbd_sdram_dat_o[30] ,
    \u_core.wbd_sdram_dat_o[29] ,
    \u_core.wbd_sdram_dat_o[28] ,
    \u_core.wbd_sdram_dat_o[27] ,
    \u_core.wbd_sdram_dat_o[26] ,
    \u_core.wbd_sdram_dat_o[25] ,
    \u_core.wbd_sdram_dat_o[24] ,
    \u_core.wbd_sdram_dat_o[23] ,
    \u_core.wbd_sdram_dat_o[22] ,
    \u_core.wbd_sdram_dat_o[21] ,
    \u_core.wbd_sdram_dat_o[20] ,
    \u_core.wbd_sdram_dat_o[19] ,
    \u_core.wbd_sdram_dat_o[18] ,
    \u_core.wbd_sdram_dat_o[17] ,
    \u_core.wbd_sdram_dat_o[16] ,
    \u_core.wbd_sdram_dat_o[15] ,
    \u_core.wbd_sdram_dat_o[14] ,
    \u_core.wbd_sdram_dat_o[13] ,
    \u_core.wbd_sdram_dat_o[12] ,
    \u_core.wbd_sdram_dat_o[11] ,
    \u_core.wbd_sdram_dat_o[10] ,
    \u_core.wbd_sdram_dat_o[9] ,
    \u_core.wbd_sdram_dat_o[8] ,
    \u_core.wbd_sdram_dat_o[7] ,
    \u_core.wbd_sdram_dat_o[6] ,
    \u_core.wbd_sdram_dat_o[5] ,
    \u_core.wbd_sdram_dat_o[4] ,
    \u_core.wbd_sdram_dat_o[3] ,
    \u_core.wbd_sdram_dat_o[2] ,
    \u_core.wbd_sdram_dat_o[1] ,
    \u_core.wbd_sdram_dat_o[0] }),
    .wb_dat_o({\u_core.wbd_sdram_dat_i[31] ,
    \u_core.wbd_sdram_dat_i[30] ,
    \u_core.wbd_sdram_dat_i[29] ,
    \u_core.wbd_sdram_dat_i[28] ,
    \u_core.wbd_sdram_dat_i[27] ,
    \u_core.wbd_sdram_dat_i[26] ,
    \u_core.wbd_sdram_dat_i[25] ,
    \u_core.wbd_sdram_dat_i[24] ,
    \u_core.wbd_sdram_dat_i[23] ,
    \u_core.wbd_sdram_dat_i[22] ,
    \u_core.wbd_sdram_dat_i[21] ,
    \u_core.wbd_sdram_dat_i[20] ,
    \u_core.wbd_sdram_dat_i[19] ,
    \u_core.wbd_sdram_dat_i[18] ,
    \u_core.wbd_sdram_dat_i[17] ,
    \u_core.wbd_sdram_dat_i[16] ,
    \u_core.wbd_sdram_dat_i[15] ,
    \u_core.wbd_sdram_dat_i[14] ,
    \u_core.wbd_sdram_dat_i[13] ,
    \u_core.wbd_sdram_dat_i[12] ,
    \u_core.wbd_sdram_dat_i[11] ,
    \u_core.wbd_sdram_dat_i[10] ,
    \u_core.wbd_sdram_dat_i[9] ,
    \u_core.wbd_sdram_dat_i[8] ,
    \u_core.wbd_sdram_dat_i[7] ,
    \u_core.wbd_sdram_dat_i[6] ,
    \u_core.wbd_sdram_dat_i[5] ,
    \u_core.wbd_sdram_dat_i[4] ,
    \u_core.wbd_sdram_dat_i[3] ,
    \u_core.wbd_sdram_dat_i[2] ,
    \u_core.wbd_sdram_dat_i[1] ,
    \u_core.wbd_sdram_dat_i[0] }),
    .wb_sel_i({\u_core.wbd_sdram_sel_o[3] ,
    \u_core.wbd_sdram_sel_o[2] ,
    \u_core.wbd_sdram_sel_o[1] ,
    \u_core.wbd_sdram_sel_o[0] }));
 spim_top \u_core.u_spi_master  (.mclk(wb_clk_i),
    .rst_n(\u_core.spi_rst_n ),
    .spi_clk(\u_core.spim_clk ),
    .spi_csn0(\u_core.spim_csn ),
    .spi_en_tx(\u_core.spi_en_tx ),
    .spi_sdi0(io_in[32]),
    .spi_sdi1(io_in[33]),
    .spi_sdi2(io_in[34]),
    .spi_sdi3(io_in[35]),
    .spi_sdo0(\u_core.spim_sdo0 ),
    .spi_sdo1(\u_core.spim_sdo1 ),
    .spi_sdo2(\u_core.spim_sdo2 ),
    .spi_sdo3(\u_core.spim_sdo3 ),
    .wbd_ack_o(\u_core.wbd_spim_ack_i ),
    .wbd_err_o(\u_core.wbd_spim_err_i ),
    .wbd_stb_i(\u_core.wbd_spim_stb_o ),
    .wbd_we_i(\u_core.wbd_spim_we_o ),
    .VPWR(vccd1),
    .VGND(vssd1),
    .events_o({_NC33,
    _NC34}),
    .spi_mode({_NC35,
    _NC36}),
    .wbd_adr_i({\u_core.wbd_spim_adr_o[31] ,
    \u_core.wbd_spim_adr_o[30] ,
    \u_core.wbd_spim_adr_o[29] ,
    \u_core.wbd_spim_adr_o[28] ,
    \u_core.wbd_spim_adr_o[27] ,
    \u_core.wbd_spim_adr_o[26] ,
    \u_core.wbd_spim_adr_o[25] ,
    \u_core.wbd_spim_adr_o[24] ,
    \u_core.wbd_spim_adr_o[23] ,
    \u_core.wbd_spim_adr_o[22] ,
    \u_core.wbd_spim_adr_o[21] ,
    \u_core.wbd_spim_adr_o[20] ,
    \u_core.wbd_spim_adr_o[19] ,
    \u_core.wbd_spim_adr_o[18] ,
    \u_core.wbd_spim_adr_o[17] ,
    \u_core.wbd_spim_adr_o[16] ,
    \u_core.wbd_spim_adr_o[15] ,
    \u_core.wbd_spim_adr_o[14] ,
    \u_core.wbd_spim_adr_o[13] ,
    \u_core.wbd_spim_adr_o[12] ,
    \u_core.wbd_spim_adr_o[11] ,
    \u_core.wbd_spim_adr_o[10] ,
    \u_core.wbd_spim_adr_o[9] ,
    \u_core.wbd_spim_adr_o[8] ,
    \u_core.wbd_spim_adr_o[7] ,
    \u_core.wbd_spim_adr_o[6] ,
    \u_core.wbd_spim_adr_o[5] ,
    \u_core.wbd_spim_adr_o[4] ,
    \u_core.wbd_spim_adr_o[3] ,
    \u_core.wbd_spim_adr_o[2] ,
    \u_core.wbd_spim_adr_o[1] ,
    \u_core.wbd_spim_adr_o[0] }),
    .wbd_dat_i({\u_core.wbd_spim_dat_o[31] ,
    \u_core.wbd_spim_dat_o[30] ,
    \u_core.wbd_spim_dat_o[29] ,
    \u_core.wbd_spim_dat_o[28] ,
    \u_core.wbd_spim_dat_o[27] ,
    \u_core.wbd_spim_dat_o[26] ,
    \u_core.wbd_spim_dat_o[25] ,
    \u_core.wbd_spim_dat_o[24] ,
    \u_core.wbd_spim_dat_o[23] ,
    \u_core.wbd_spim_dat_o[22] ,
    \u_core.wbd_spim_dat_o[21] ,
    \u_core.wbd_spim_dat_o[20] ,
    \u_core.wbd_spim_dat_o[19] ,
    \u_core.wbd_spim_dat_o[18] ,
    \u_core.wbd_spim_dat_o[17] ,
    \u_core.wbd_spim_dat_o[16] ,
    \u_core.wbd_spim_dat_o[15] ,
    \u_core.wbd_spim_dat_o[14] ,
    \u_core.wbd_spim_dat_o[13] ,
    \u_core.wbd_spim_dat_o[12] ,
    \u_core.wbd_spim_dat_o[11] ,
    \u_core.wbd_spim_dat_o[10] ,
    \u_core.wbd_spim_dat_o[9] ,
    \u_core.wbd_spim_dat_o[8] ,
    \u_core.wbd_spim_dat_o[7] ,
    \u_core.wbd_spim_dat_o[6] ,
    \u_core.wbd_spim_dat_o[5] ,
    \u_core.wbd_spim_dat_o[4] ,
    \u_core.wbd_spim_dat_o[3] ,
    \u_core.wbd_spim_dat_o[2] ,
    \u_core.wbd_spim_dat_o[1] ,
    \u_core.wbd_spim_dat_o[0] }),
    .wbd_dat_o({\u_core.wbd_spim_dat_i[31] ,
    \u_core.wbd_spim_dat_i[30] ,
    \u_core.wbd_spim_dat_i[29] ,
    \u_core.wbd_spim_dat_i[28] ,
    \u_core.wbd_spim_dat_i[27] ,
    \u_core.wbd_spim_dat_i[26] ,
    \u_core.wbd_spim_dat_i[25] ,
    \u_core.wbd_spim_dat_i[24] ,
    \u_core.wbd_spim_dat_i[23] ,
    \u_core.wbd_spim_dat_i[22] ,
    \u_core.wbd_spim_dat_i[21] ,
    \u_core.wbd_spim_dat_i[20] ,
    \u_core.wbd_spim_dat_i[19] ,
    \u_core.wbd_spim_dat_i[18] ,
    \u_core.wbd_spim_dat_i[17] ,
    \u_core.wbd_spim_dat_i[16] ,
    \u_core.wbd_spim_dat_i[15] ,
    \u_core.wbd_spim_dat_i[14] ,
    \u_core.wbd_spim_dat_i[13] ,
    \u_core.wbd_spim_dat_i[12] ,
    \u_core.wbd_spim_dat_i[11] ,
    \u_core.wbd_spim_dat_i[10] ,
    \u_core.wbd_spim_dat_i[9] ,
    \u_core.wbd_spim_dat_i[8] ,
    \u_core.wbd_spim_dat_i[7] ,
    \u_core.wbd_spim_dat_i[6] ,
    \u_core.wbd_spim_dat_i[5] ,
    \u_core.wbd_spim_dat_i[4] ,
    \u_core.wbd_spim_dat_i[3] ,
    \u_core.wbd_spim_dat_i[2] ,
    \u_core.wbd_spim_dat_i[1] ,
    \u_core.wbd_spim_dat_i[0] }),
    .wbd_sel_i({\u_core.wbd_spim_sel_o[3] ,
    \u_core.wbd_spim_sel_o[2] ,
    \u_core.wbd_spim_sel_o[1] ,
    \u_core.wbd_spim_sel_o[0] }));
endmodule
