module user_project_wrapper (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    vccd1,
    vssd1,
    analog_io,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input vccd1;
 input vssd1;
 inout [28:0] analog_io;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 glbl_cfg u_glbl_cfg (.cfg_sdr_en(cfg_sdr_en),
    .mclk(wbd_clk_glbl),
    .reg_ack(wbd_glbl_ack_i),
    .reg_cs(wbd_glbl_stb_o),
    .reg_wr(wbd_glbl_we_o),
    .reset_n(wbd_int_rst_n),
    .sdr_init_done(sdr_init_done),
    .soft_irq(soft_irq),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .cfg_colbits({\cfg_colbits[1] ,
    \cfg_colbits[0] }),
    .cfg_req_depth({\cfg_req_depth[1] ,
    \cfg_req_depth[0] }),
    .cfg_sdr_cas({\cfg_sdr_cas[2] ,
    \cfg_sdr_cas[1] ,
    \cfg_sdr_cas[0] }),
    .cfg_sdr_mode_reg({\cfg_sdr_mode_reg[12] ,
    \cfg_sdr_mode_reg[11] ,
    \cfg_sdr_mode_reg[10] ,
    \cfg_sdr_mode_reg[9] ,
    \cfg_sdr_mode_reg[8] ,
    \cfg_sdr_mode_reg[7] ,
    \cfg_sdr_mode_reg[6] ,
    \cfg_sdr_mode_reg[5] ,
    \cfg_sdr_mode_reg[4] ,
    \cfg_sdr_mode_reg[3] ,
    \cfg_sdr_mode_reg[2] ,
    \cfg_sdr_mode_reg[1] ,
    \cfg_sdr_mode_reg[0] }),
    .cfg_sdr_rfmax({\cfg_sdr_rfmax[2] ,
    \cfg_sdr_rfmax[1] ,
    \cfg_sdr_rfmax[0] }),
    .cfg_sdr_rfsh({\cfg_sdr_rfsh[11] ,
    \cfg_sdr_rfsh[10] ,
    \cfg_sdr_rfsh[9] ,
    \cfg_sdr_rfsh[8] ,
    \cfg_sdr_rfsh[7] ,
    \cfg_sdr_rfsh[6] ,
    \cfg_sdr_rfsh[5] ,
    \cfg_sdr_rfsh[4] ,
    \cfg_sdr_rfsh[3] ,
    \cfg_sdr_rfsh[2] ,
    \cfg_sdr_rfsh[1] ,
    \cfg_sdr_rfsh[0] }),
    .cfg_sdr_tras_d({\cfg_sdr_tras_d[3] ,
    \cfg_sdr_tras_d[2] ,
    \cfg_sdr_tras_d[1] ,
    \cfg_sdr_tras_d[0] }),
    .cfg_sdr_trcar_d({\cfg_sdr_trcar_d[3] ,
    \cfg_sdr_trcar_d[2] ,
    \cfg_sdr_trcar_d[1] ,
    \cfg_sdr_trcar_d[0] }),
    .cfg_sdr_trcd_d({\cfg_sdr_trcd_d[3] ,
    \cfg_sdr_trcd_d[2] ,
    \cfg_sdr_trcd_d[1] ,
    \cfg_sdr_trcd_d[0] }),
    .cfg_sdr_trp_d({\cfg_sdr_trp_d[3] ,
    \cfg_sdr_trp_d[2] ,
    \cfg_sdr_trp_d[1] ,
    \cfg_sdr_trp_d[0] }),
    .cfg_sdr_twr_d({\cfg_sdr_twr_d[3] ,
    \cfg_sdr_twr_d[2] ,
    \cfg_sdr_twr_d[1] ,
    \cfg_sdr_twr_d[0] }),
    .cfg_sdr_width({\cfg_sdr_width[1] ,
    \cfg_sdr_width[0] }),
    .fuse_mhartid({\fuse_mhartid[31] ,
    \fuse_mhartid[30] ,
    \fuse_mhartid[29] ,
    \fuse_mhartid[28] ,
    \fuse_mhartid[27] ,
    \fuse_mhartid[26] ,
    \fuse_mhartid[25] ,
    \fuse_mhartid[24] ,
    \fuse_mhartid[23] ,
    \fuse_mhartid[22] ,
    \fuse_mhartid[21] ,
    \fuse_mhartid[20] ,
    \fuse_mhartid[19] ,
    \fuse_mhartid[18] ,
    \fuse_mhartid[17] ,
    \fuse_mhartid[16] ,
    \fuse_mhartid[15] ,
    \fuse_mhartid[14] ,
    \fuse_mhartid[13] ,
    \fuse_mhartid[12] ,
    \fuse_mhartid[11] ,
    \fuse_mhartid[10] ,
    \fuse_mhartid[9] ,
    \fuse_mhartid[8] ,
    \fuse_mhartid[7] ,
    \fuse_mhartid[6] ,
    \fuse_mhartid[5] ,
    \fuse_mhartid[4] ,
    \fuse_mhartid[3] ,
    \fuse_mhartid[2] ,
    \fuse_mhartid[1] ,
    \fuse_mhartid[0] }),
    .irq_lines({\irq_lines[15] ,
    \irq_lines[14] ,
    \irq_lines[13] ,
    \irq_lines[12] ,
    \irq_lines[11] ,
    \irq_lines[10] ,
    \irq_lines[9] ,
    \irq_lines[8] ,
    \irq_lines[7] ,
    \irq_lines[6] ,
    \irq_lines[5] ,
    \irq_lines[4] ,
    \irq_lines[3] ,
    \irq_lines[2] ,
    \irq_lines[1] ,
    \irq_lines[0] }),
    .reg_addr({\wbd_glbl_adr_o[7] ,
    \wbd_glbl_adr_o[6] ,
    \wbd_glbl_adr_o[5] ,
    \wbd_glbl_adr_o[4] ,
    \wbd_glbl_adr_o[3] ,
    \wbd_glbl_adr_o[2] ,
    \wbd_glbl_adr_o[1] ,
    \wbd_glbl_adr_o[0] }),
    .reg_be({\wbd_glbl_sel_o[3] ,
    \wbd_glbl_sel_o[2] ,
    \wbd_glbl_sel_o[1] ,
    \wbd_glbl_sel_o[0] }),
    .reg_rdata({\wbd_glbl_dat_i[31] ,
    \wbd_glbl_dat_i[30] ,
    \wbd_glbl_dat_i[29] ,
    \wbd_glbl_dat_i[28] ,
    \wbd_glbl_dat_i[27] ,
    \wbd_glbl_dat_i[26] ,
    \wbd_glbl_dat_i[25] ,
    \wbd_glbl_dat_i[24] ,
    \wbd_glbl_dat_i[23] ,
    \wbd_glbl_dat_i[22] ,
    \wbd_glbl_dat_i[21] ,
    \wbd_glbl_dat_i[20] ,
    \wbd_glbl_dat_i[19] ,
    \wbd_glbl_dat_i[18] ,
    \wbd_glbl_dat_i[17] ,
    \wbd_glbl_dat_i[16] ,
    \wbd_glbl_dat_i[15] ,
    \wbd_glbl_dat_i[14] ,
    \wbd_glbl_dat_i[13] ,
    \wbd_glbl_dat_i[12] ,
    \wbd_glbl_dat_i[11] ,
    \wbd_glbl_dat_i[10] ,
    \wbd_glbl_dat_i[9] ,
    \wbd_glbl_dat_i[8] ,
    \wbd_glbl_dat_i[7] ,
    \wbd_glbl_dat_i[6] ,
    \wbd_glbl_dat_i[5] ,
    \wbd_glbl_dat_i[4] ,
    \wbd_glbl_dat_i[3] ,
    \wbd_glbl_dat_i[2] ,
    \wbd_glbl_dat_i[1] ,
    \wbd_glbl_dat_i[0] }),
    .reg_wdata({\wbd_glbl_dat_o[31] ,
    \wbd_glbl_dat_o[30] ,
    \wbd_glbl_dat_o[29] ,
    \wbd_glbl_dat_o[28] ,
    \wbd_glbl_dat_o[27] ,
    \wbd_glbl_dat_o[26] ,
    \wbd_glbl_dat_o[25] ,
    \wbd_glbl_dat_o[24] ,
    \wbd_glbl_dat_o[23] ,
    \wbd_glbl_dat_o[22] ,
    \wbd_glbl_dat_o[21] ,
    \wbd_glbl_dat_o[20] ,
    \wbd_glbl_dat_o[19] ,
    \wbd_glbl_dat_o[18] ,
    \wbd_glbl_dat_o[17] ,
    \wbd_glbl_dat_o[16] ,
    \wbd_glbl_dat_o[15] ,
    \wbd_glbl_dat_o[14] ,
    \wbd_glbl_dat_o[13] ,
    \wbd_glbl_dat_o[12] ,
    \wbd_glbl_dat_o[11] ,
    \wbd_glbl_dat_o[10] ,
    \wbd_glbl_dat_o[9] ,
    \wbd_glbl_dat_o[8] ,
    \wbd_glbl_dat_o[7] ,
    \wbd_glbl_dat_o[6] ,
    \wbd_glbl_dat_o[5] ,
    \wbd_glbl_dat_o[4] ,
    \wbd_glbl_dat_o[3] ,
    \wbd_glbl_dat_o[2] ,
    \wbd_glbl_dat_o[1] ,
    \wbd_glbl_dat_o[0] }),
    .user_irq({user_irq[2],
    user_irq[1],
    user_irq[0]}));
 wb_interconnect u_intercon (.clk_i(wbd_clk_wi),
    .m0_wbd_ack_o(wbd_int_ack_o),
    .m0_wbd_cyc_i(wbd_int_cyc_i),
    .m0_wbd_err_o(wbd_int_err_o),
    .m0_wbd_stb_i(wbd_int_stb_i),
    .m0_wbd_we_i(wbd_int_we_i),
    .m1_wbd_ack_o(wbd_riscv_imem_ack_o),
    .m1_wbd_cyc_i(wbd_riscv_imem_stb_i),
    .m1_wbd_err_o(wbd_riscv_imem_err_o),
    .m1_wbd_stb_i(wbd_riscv_imem_stb_i),
    .m1_wbd_we_i(wbd_riscv_imem_we_i),
    .m2_wbd_ack_o(wbd_riscv_dmem_ack_o),
    .m2_wbd_cyc_i(wbd_riscv_dmem_stb_i),
    .m2_wbd_err_o(wbd_riscv_dmem_err_o),
    .m2_wbd_stb_i(wbd_riscv_dmem_stb_i),
    .m2_wbd_we_i(wbd_riscv_dmem_we_i),
    .rst_n(wbd_int_rst_n),
    .s0_wbd_ack_i(wbd_spim_ack_i),
    .s0_wbd_cyc_o(wbd_spim_cyc_o),
    .s0_wbd_stb_o(wbd_spim_stb_o),
    .s0_wbd_we_o(wbd_spim_we_o),
    .s1_wbd_ack_i(wbd_sdram_ack_i),
    .s1_wbd_cyc_o(wbd_sdram_cyc_o),
    .s1_wbd_stb_o(wbd_sdram_stb_o),
    .s1_wbd_we_o(wbd_sdram_we_o),
    .s2_wbd_ack_i(wbd_glbl_ack_i),
    .s2_wbd_cyc_o(wbd_glbl_cyc_o),
    .s2_wbd_stb_o(wbd_glbl_stb_o),
    .s2_wbd_we_o(wbd_glbl_we_o),
    .s3_wbd_ack_i(wbd_uart_ack_i),
    .s3_wbd_cyc_o(wbd_uart_cyc_o),
    .s3_wbd_sel_o(wbd_uart_sel_o),
    .s3_wbd_stb_o(wbd_uart_stb_o),
    .s3_wbd_we_o(wbd_uart_we_o),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .m0_wbd_adr_i({\wbd_int_adr_i[31] ,
    \wbd_int_adr_i[30] ,
    \wbd_int_adr_i[29] ,
    \wbd_int_adr_i[28] ,
    \wbd_int_adr_i[27] ,
    \wbd_int_adr_i[26] ,
    \wbd_int_adr_i[25] ,
    \wbd_int_adr_i[24] ,
    \wbd_int_adr_i[23] ,
    \wbd_int_adr_i[22] ,
    \wbd_int_adr_i[21] ,
    \wbd_int_adr_i[20] ,
    \wbd_int_adr_i[19] ,
    \wbd_int_adr_i[18] ,
    \wbd_int_adr_i[17] ,
    \wbd_int_adr_i[16] ,
    \wbd_int_adr_i[15] ,
    \wbd_int_adr_i[14] ,
    \wbd_int_adr_i[13] ,
    \wbd_int_adr_i[12] ,
    \wbd_int_adr_i[11] ,
    \wbd_int_adr_i[10] ,
    \wbd_int_adr_i[9] ,
    \wbd_int_adr_i[8] ,
    \wbd_int_adr_i[7] ,
    \wbd_int_adr_i[6] ,
    \wbd_int_adr_i[5] ,
    \wbd_int_adr_i[4] ,
    \wbd_int_adr_i[3] ,
    \wbd_int_adr_i[2] ,
    \wbd_int_adr_i[1] ,
    \wbd_int_adr_i[0] }),
    .m0_wbd_dat_i({\wbd_int_dat_i[31] ,
    \wbd_int_dat_i[30] ,
    \wbd_int_dat_i[29] ,
    \wbd_int_dat_i[28] ,
    \wbd_int_dat_i[27] ,
    \wbd_int_dat_i[26] ,
    \wbd_int_dat_i[25] ,
    \wbd_int_dat_i[24] ,
    \wbd_int_dat_i[23] ,
    \wbd_int_dat_i[22] ,
    \wbd_int_dat_i[21] ,
    \wbd_int_dat_i[20] ,
    \wbd_int_dat_i[19] ,
    \wbd_int_dat_i[18] ,
    \wbd_int_dat_i[17] ,
    \wbd_int_dat_i[16] ,
    \wbd_int_dat_i[15] ,
    \wbd_int_dat_i[14] ,
    \wbd_int_dat_i[13] ,
    \wbd_int_dat_i[12] ,
    \wbd_int_dat_i[11] ,
    \wbd_int_dat_i[10] ,
    \wbd_int_dat_i[9] ,
    \wbd_int_dat_i[8] ,
    \wbd_int_dat_i[7] ,
    \wbd_int_dat_i[6] ,
    \wbd_int_dat_i[5] ,
    \wbd_int_dat_i[4] ,
    \wbd_int_dat_i[3] ,
    \wbd_int_dat_i[2] ,
    \wbd_int_dat_i[1] ,
    \wbd_int_dat_i[0] }),
    .m0_wbd_dat_o({\wbd_int_dat_o[31] ,
    \wbd_int_dat_o[30] ,
    \wbd_int_dat_o[29] ,
    \wbd_int_dat_o[28] ,
    \wbd_int_dat_o[27] ,
    \wbd_int_dat_o[26] ,
    \wbd_int_dat_o[25] ,
    \wbd_int_dat_o[24] ,
    \wbd_int_dat_o[23] ,
    \wbd_int_dat_o[22] ,
    \wbd_int_dat_o[21] ,
    \wbd_int_dat_o[20] ,
    \wbd_int_dat_o[19] ,
    \wbd_int_dat_o[18] ,
    \wbd_int_dat_o[17] ,
    \wbd_int_dat_o[16] ,
    \wbd_int_dat_o[15] ,
    \wbd_int_dat_o[14] ,
    \wbd_int_dat_o[13] ,
    \wbd_int_dat_o[12] ,
    \wbd_int_dat_o[11] ,
    \wbd_int_dat_o[10] ,
    \wbd_int_dat_o[9] ,
    \wbd_int_dat_o[8] ,
    \wbd_int_dat_o[7] ,
    \wbd_int_dat_o[6] ,
    \wbd_int_dat_o[5] ,
    \wbd_int_dat_o[4] ,
    \wbd_int_dat_o[3] ,
    \wbd_int_dat_o[2] ,
    \wbd_int_dat_o[1] ,
    \wbd_int_dat_o[0] }),
    .m0_wbd_sel_i({\wbd_int_sel_i[3] ,
    \wbd_int_sel_i[2] ,
    \wbd_int_sel_i[1] ,
    \wbd_int_sel_i[0] }),
    .m1_wbd_adr_i({\wbd_riscv_imem_adr_i[31] ,
    \wbd_riscv_imem_adr_i[30] ,
    \wbd_riscv_imem_adr_i[29] ,
    \wbd_riscv_imem_adr_i[28] ,
    \wbd_riscv_imem_adr_i[27] ,
    \wbd_riscv_imem_adr_i[26] ,
    \wbd_riscv_imem_adr_i[25] ,
    \wbd_riscv_imem_adr_i[24] ,
    \wbd_riscv_imem_adr_i[23] ,
    \wbd_riscv_imem_adr_i[22] ,
    \wbd_riscv_imem_adr_i[21] ,
    \wbd_riscv_imem_adr_i[20] ,
    \wbd_riscv_imem_adr_i[19] ,
    \wbd_riscv_imem_adr_i[18] ,
    \wbd_riscv_imem_adr_i[17] ,
    \wbd_riscv_imem_adr_i[16] ,
    \wbd_riscv_imem_adr_i[15] ,
    \wbd_riscv_imem_adr_i[14] ,
    \wbd_riscv_imem_adr_i[13] ,
    \wbd_riscv_imem_adr_i[12] ,
    \wbd_riscv_imem_adr_i[11] ,
    \wbd_riscv_imem_adr_i[10] ,
    \wbd_riscv_imem_adr_i[9] ,
    \wbd_riscv_imem_adr_i[8] ,
    \wbd_riscv_imem_adr_i[7] ,
    \wbd_riscv_imem_adr_i[6] ,
    \wbd_riscv_imem_adr_i[5] ,
    \wbd_riscv_imem_adr_i[4] ,
    \wbd_riscv_imem_adr_i[3] ,
    \wbd_riscv_imem_adr_i[2] ,
    \wbd_riscv_imem_adr_i[1] ,
    \wbd_riscv_imem_adr_i[0] }),
    .m1_wbd_dat_i({\wbd_riscv_imem_dat_i[31] ,
    \wbd_riscv_imem_dat_i[30] ,
    \wbd_riscv_imem_dat_i[29] ,
    \wbd_riscv_imem_dat_i[28] ,
    \wbd_riscv_imem_dat_i[27] ,
    \wbd_riscv_imem_dat_i[26] ,
    \wbd_riscv_imem_dat_i[25] ,
    \wbd_riscv_imem_dat_i[24] ,
    \wbd_riscv_imem_dat_i[23] ,
    \wbd_riscv_imem_dat_i[22] ,
    \wbd_riscv_imem_dat_i[21] ,
    \wbd_riscv_imem_dat_i[20] ,
    \wbd_riscv_imem_dat_i[19] ,
    \wbd_riscv_imem_dat_i[18] ,
    \wbd_riscv_imem_dat_i[17] ,
    \wbd_riscv_imem_dat_i[16] ,
    \wbd_riscv_imem_dat_i[15] ,
    \wbd_riscv_imem_dat_i[14] ,
    \wbd_riscv_imem_dat_i[13] ,
    \wbd_riscv_imem_dat_i[12] ,
    \wbd_riscv_imem_dat_i[11] ,
    \wbd_riscv_imem_dat_i[10] ,
    \wbd_riscv_imem_dat_i[9] ,
    \wbd_riscv_imem_dat_i[8] ,
    \wbd_riscv_imem_dat_i[7] ,
    \wbd_riscv_imem_dat_i[6] ,
    \wbd_riscv_imem_dat_i[5] ,
    \wbd_riscv_imem_dat_i[4] ,
    \wbd_riscv_imem_dat_i[3] ,
    \wbd_riscv_imem_dat_i[2] ,
    \wbd_riscv_imem_dat_i[1] ,
    \wbd_riscv_imem_dat_i[0] }),
    .m1_wbd_dat_o({\wbd_riscv_imem_dat_o[31] ,
    \wbd_riscv_imem_dat_o[30] ,
    \wbd_riscv_imem_dat_o[29] ,
    \wbd_riscv_imem_dat_o[28] ,
    \wbd_riscv_imem_dat_o[27] ,
    \wbd_riscv_imem_dat_o[26] ,
    \wbd_riscv_imem_dat_o[25] ,
    \wbd_riscv_imem_dat_o[24] ,
    \wbd_riscv_imem_dat_o[23] ,
    \wbd_riscv_imem_dat_o[22] ,
    \wbd_riscv_imem_dat_o[21] ,
    \wbd_riscv_imem_dat_o[20] ,
    \wbd_riscv_imem_dat_o[19] ,
    \wbd_riscv_imem_dat_o[18] ,
    \wbd_riscv_imem_dat_o[17] ,
    \wbd_riscv_imem_dat_o[16] ,
    \wbd_riscv_imem_dat_o[15] ,
    \wbd_riscv_imem_dat_o[14] ,
    \wbd_riscv_imem_dat_o[13] ,
    \wbd_riscv_imem_dat_o[12] ,
    \wbd_riscv_imem_dat_o[11] ,
    \wbd_riscv_imem_dat_o[10] ,
    \wbd_riscv_imem_dat_o[9] ,
    \wbd_riscv_imem_dat_o[8] ,
    \wbd_riscv_imem_dat_o[7] ,
    \wbd_riscv_imem_dat_o[6] ,
    \wbd_riscv_imem_dat_o[5] ,
    \wbd_riscv_imem_dat_o[4] ,
    \wbd_riscv_imem_dat_o[3] ,
    \wbd_riscv_imem_dat_o[2] ,
    \wbd_riscv_imem_dat_o[1] ,
    \wbd_riscv_imem_dat_o[0] }),
    .m1_wbd_sel_i({\wbd_riscv_imem_sel_i[3] ,
    \wbd_riscv_imem_sel_i[2] ,
    \wbd_riscv_imem_sel_i[1] ,
    \wbd_riscv_imem_sel_i[0] }),
    .m2_wbd_adr_i({\wbd_riscv_dmem_adr_i[31] ,
    \wbd_riscv_dmem_adr_i[30] ,
    \wbd_riscv_dmem_adr_i[29] ,
    \wbd_riscv_dmem_adr_i[28] ,
    \wbd_riscv_dmem_adr_i[27] ,
    \wbd_riscv_dmem_adr_i[26] ,
    \wbd_riscv_dmem_adr_i[25] ,
    \wbd_riscv_dmem_adr_i[24] ,
    \wbd_riscv_dmem_adr_i[23] ,
    \wbd_riscv_dmem_adr_i[22] ,
    \wbd_riscv_dmem_adr_i[21] ,
    \wbd_riscv_dmem_adr_i[20] ,
    \wbd_riscv_dmem_adr_i[19] ,
    \wbd_riscv_dmem_adr_i[18] ,
    \wbd_riscv_dmem_adr_i[17] ,
    \wbd_riscv_dmem_adr_i[16] ,
    \wbd_riscv_dmem_adr_i[15] ,
    \wbd_riscv_dmem_adr_i[14] ,
    \wbd_riscv_dmem_adr_i[13] ,
    \wbd_riscv_dmem_adr_i[12] ,
    \wbd_riscv_dmem_adr_i[11] ,
    \wbd_riscv_dmem_adr_i[10] ,
    \wbd_riscv_dmem_adr_i[9] ,
    \wbd_riscv_dmem_adr_i[8] ,
    \wbd_riscv_dmem_adr_i[7] ,
    \wbd_riscv_dmem_adr_i[6] ,
    \wbd_riscv_dmem_adr_i[5] ,
    \wbd_riscv_dmem_adr_i[4] ,
    \wbd_riscv_dmem_adr_i[3] ,
    \wbd_riscv_dmem_adr_i[2] ,
    \wbd_riscv_dmem_adr_i[1] ,
    \wbd_riscv_dmem_adr_i[0] }),
    .m2_wbd_dat_i({\wbd_riscv_dmem_dat_i[31] ,
    \wbd_riscv_dmem_dat_i[30] ,
    \wbd_riscv_dmem_dat_i[29] ,
    \wbd_riscv_dmem_dat_i[28] ,
    \wbd_riscv_dmem_dat_i[27] ,
    \wbd_riscv_dmem_dat_i[26] ,
    \wbd_riscv_dmem_dat_i[25] ,
    \wbd_riscv_dmem_dat_i[24] ,
    \wbd_riscv_dmem_dat_i[23] ,
    \wbd_riscv_dmem_dat_i[22] ,
    \wbd_riscv_dmem_dat_i[21] ,
    \wbd_riscv_dmem_dat_i[20] ,
    \wbd_riscv_dmem_dat_i[19] ,
    \wbd_riscv_dmem_dat_i[18] ,
    \wbd_riscv_dmem_dat_i[17] ,
    \wbd_riscv_dmem_dat_i[16] ,
    \wbd_riscv_dmem_dat_i[15] ,
    \wbd_riscv_dmem_dat_i[14] ,
    \wbd_riscv_dmem_dat_i[13] ,
    \wbd_riscv_dmem_dat_i[12] ,
    \wbd_riscv_dmem_dat_i[11] ,
    \wbd_riscv_dmem_dat_i[10] ,
    \wbd_riscv_dmem_dat_i[9] ,
    \wbd_riscv_dmem_dat_i[8] ,
    \wbd_riscv_dmem_dat_i[7] ,
    \wbd_riscv_dmem_dat_i[6] ,
    \wbd_riscv_dmem_dat_i[5] ,
    \wbd_riscv_dmem_dat_i[4] ,
    \wbd_riscv_dmem_dat_i[3] ,
    \wbd_riscv_dmem_dat_i[2] ,
    \wbd_riscv_dmem_dat_i[1] ,
    \wbd_riscv_dmem_dat_i[0] }),
    .m2_wbd_dat_o({\wbd_riscv_dmem_dat_o[31] ,
    \wbd_riscv_dmem_dat_o[30] ,
    \wbd_riscv_dmem_dat_o[29] ,
    \wbd_riscv_dmem_dat_o[28] ,
    \wbd_riscv_dmem_dat_o[27] ,
    \wbd_riscv_dmem_dat_o[26] ,
    \wbd_riscv_dmem_dat_o[25] ,
    \wbd_riscv_dmem_dat_o[24] ,
    \wbd_riscv_dmem_dat_o[23] ,
    \wbd_riscv_dmem_dat_o[22] ,
    \wbd_riscv_dmem_dat_o[21] ,
    \wbd_riscv_dmem_dat_o[20] ,
    \wbd_riscv_dmem_dat_o[19] ,
    \wbd_riscv_dmem_dat_o[18] ,
    \wbd_riscv_dmem_dat_o[17] ,
    \wbd_riscv_dmem_dat_o[16] ,
    \wbd_riscv_dmem_dat_o[15] ,
    \wbd_riscv_dmem_dat_o[14] ,
    \wbd_riscv_dmem_dat_o[13] ,
    \wbd_riscv_dmem_dat_o[12] ,
    \wbd_riscv_dmem_dat_o[11] ,
    \wbd_riscv_dmem_dat_o[10] ,
    \wbd_riscv_dmem_dat_o[9] ,
    \wbd_riscv_dmem_dat_o[8] ,
    \wbd_riscv_dmem_dat_o[7] ,
    \wbd_riscv_dmem_dat_o[6] ,
    \wbd_riscv_dmem_dat_o[5] ,
    \wbd_riscv_dmem_dat_o[4] ,
    \wbd_riscv_dmem_dat_o[3] ,
    \wbd_riscv_dmem_dat_o[2] ,
    \wbd_riscv_dmem_dat_o[1] ,
    \wbd_riscv_dmem_dat_o[0] }),
    .m2_wbd_sel_i({\wbd_riscv_dmem_sel_i[3] ,
    \wbd_riscv_dmem_sel_i[2] ,
    \wbd_riscv_dmem_sel_i[1] ,
    \wbd_riscv_dmem_sel_i[0] }),
    .s0_wbd_adr_o({\wbd_spim_adr_o[31] ,
    \wbd_spim_adr_o[30] ,
    \wbd_spim_adr_o[29] ,
    \wbd_spim_adr_o[28] ,
    \wbd_spim_adr_o[27] ,
    \wbd_spim_adr_o[26] ,
    \wbd_spim_adr_o[25] ,
    \wbd_spim_adr_o[24] ,
    \wbd_spim_adr_o[23] ,
    \wbd_spim_adr_o[22] ,
    \wbd_spim_adr_o[21] ,
    \wbd_spim_adr_o[20] ,
    \wbd_spim_adr_o[19] ,
    \wbd_spim_adr_o[18] ,
    \wbd_spim_adr_o[17] ,
    \wbd_spim_adr_o[16] ,
    \wbd_spim_adr_o[15] ,
    \wbd_spim_adr_o[14] ,
    \wbd_spim_adr_o[13] ,
    \wbd_spim_adr_o[12] ,
    \wbd_spim_adr_o[11] ,
    \wbd_spim_adr_o[10] ,
    \wbd_spim_adr_o[9] ,
    \wbd_spim_adr_o[8] ,
    \wbd_spim_adr_o[7] ,
    \wbd_spim_adr_o[6] ,
    \wbd_spim_adr_o[5] ,
    \wbd_spim_adr_o[4] ,
    \wbd_spim_adr_o[3] ,
    \wbd_spim_adr_o[2] ,
    \wbd_spim_adr_o[1] ,
    \wbd_spim_adr_o[0] }),
    .s0_wbd_dat_i({\wbd_spim_dat_i[31] ,
    \wbd_spim_dat_i[30] ,
    \wbd_spim_dat_i[29] ,
    \wbd_spim_dat_i[28] ,
    \wbd_spim_dat_i[27] ,
    \wbd_spim_dat_i[26] ,
    \wbd_spim_dat_i[25] ,
    \wbd_spim_dat_i[24] ,
    \wbd_spim_dat_i[23] ,
    \wbd_spim_dat_i[22] ,
    \wbd_spim_dat_i[21] ,
    \wbd_spim_dat_i[20] ,
    \wbd_spim_dat_i[19] ,
    \wbd_spim_dat_i[18] ,
    \wbd_spim_dat_i[17] ,
    \wbd_spim_dat_i[16] ,
    \wbd_spim_dat_i[15] ,
    \wbd_spim_dat_i[14] ,
    \wbd_spim_dat_i[13] ,
    \wbd_spim_dat_i[12] ,
    \wbd_spim_dat_i[11] ,
    \wbd_spim_dat_i[10] ,
    \wbd_spim_dat_i[9] ,
    \wbd_spim_dat_i[8] ,
    \wbd_spim_dat_i[7] ,
    \wbd_spim_dat_i[6] ,
    \wbd_spim_dat_i[5] ,
    \wbd_spim_dat_i[4] ,
    \wbd_spim_dat_i[3] ,
    \wbd_spim_dat_i[2] ,
    \wbd_spim_dat_i[1] ,
    \wbd_spim_dat_i[0] }),
    .s0_wbd_dat_o({\wbd_spim_dat_o[31] ,
    \wbd_spim_dat_o[30] ,
    \wbd_spim_dat_o[29] ,
    \wbd_spim_dat_o[28] ,
    \wbd_spim_dat_o[27] ,
    \wbd_spim_dat_o[26] ,
    \wbd_spim_dat_o[25] ,
    \wbd_spim_dat_o[24] ,
    \wbd_spim_dat_o[23] ,
    \wbd_spim_dat_o[22] ,
    \wbd_spim_dat_o[21] ,
    \wbd_spim_dat_o[20] ,
    \wbd_spim_dat_o[19] ,
    \wbd_spim_dat_o[18] ,
    \wbd_spim_dat_o[17] ,
    \wbd_spim_dat_o[16] ,
    \wbd_spim_dat_o[15] ,
    \wbd_spim_dat_o[14] ,
    \wbd_spim_dat_o[13] ,
    \wbd_spim_dat_o[12] ,
    \wbd_spim_dat_o[11] ,
    \wbd_spim_dat_o[10] ,
    \wbd_spim_dat_o[9] ,
    \wbd_spim_dat_o[8] ,
    \wbd_spim_dat_o[7] ,
    \wbd_spim_dat_o[6] ,
    \wbd_spim_dat_o[5] ,
    \wbd_spim_dat_o[4] ,
    \wbd_spim_dat_o[3] ,
    \wbd_spim_dat_o[2] ,
    \wbd_spim_dat_o[1] ,
    \wbd_spim_dat_o[0] }),
    .s0_wbd_sel_o({\wbd_spim_sel_o[3] ,
    \wbd_spim_sel_o[2] ,
    \wbd_spim_sel_o[1] ,
    \wbd_spim_sel_o[0] }),
    .s1_wbd_adr_o({\wbd_sdram_adr_o[31] ,
    \wbd_sdram_adr_o[30] ,
    \wbd_sdram_adr_o[29] ,
    \wbd_sdram_adr_o[28] ,
    \wbd_sdram_adr_o[27] ,
    \wbd_sdram_adr_o[26] ,
    \wbd_sdram_adr_o[25] ,
    \wbd_sdram_adr_o[24] ,
    \wbd_sdram_adr_o[23] ,
    \wbd_sdram_adr_o[22] ,
    \wbd_sdram_adr_o[21] ,
    \wbd_sdram_adr_o[20] ,
    \wbd_sdram_adr_o[19] ,
    \wbd_sdram_adr_o[18] ,
    \wbd_sdram_adr_o[17] ,
    \wbd_sdram_adr_o[16] ,
    \wbd_sdram_adr_o[15] ,
    \wbd_sdram_adr_o[14] ,
    \wbd_sdram_adr_o[13] ,
    \wbd_sdram_adr_o[12] ,
    \wbd_sdram_adr_o[11] ,
    \wbd_sdram_adr_o[10] ,
    \wbd_sdram_adr_o[9] ,
    \wbd_sdram_adr_o[8] ,
    \wbd_sdram_adr_o[7] ,
    \wbd_sdram_adr_o[6] ,
    \wbd_sdram_adr_o[5] ,
    \wbd_sdram_adr_o[4] ,
    \wbd_sdram_adr_o[3] ,
    \wbd_sdram_adr_o[2] ,
    \wbd_sdram_adr_o[1] ,
    \wbd_sdram_adr_o[0] }),
    .s1_wbd_dat_i({\wbd_sdram_dat_i[31] ,
    \wbd_sdram_dat_i[30] ,
    \wbd_sdram_dat_i[29] ,
    \wbd_sdram_dat_i[28] ,
    \wbd_sdram_dat_i[27] ,
    \wbd_sdram_dat_i[26] ,
    \wbd_sdram_dat_i[25] ,
    \wbd_sdram_dat_i[24] ,
    \wbd_sdram_dat_i[23] ,
    \wbd_sdram_dat_i[22] ,
    \wbd_sdram_dat_i[21] ,
    \wbd_sdram_dat_i[20] ,
    \wbd_sdram_dat_i[19] ,
    \wbd_sdram_dat_i[18] ,
    \wbd_sdram_dat_i[17] ,
    \wbd_sdram_dat_i[16] ,
    \wbd_sdram_dat_i[15] ,
    \wbd_sdram_dat_i[14] ,
    \wbd_sdram_dat_i[13] ,
    \wbd_sdram_dat_i[12] ,
    \wbd_sdram_dat_i[11] ,
    \wbd_sdram_dat_i[10] ,
    \wbd_sdram_dat_i[9] ,
    \wbd_sdram_dat_i[8] ,
    \wbd_sdram_dat_i[7] ,
    \wbd_sdram_dat_i[6] ,
    \wbd_sdram_dat_i[5] ,
    \wbd_sdram_dat_i[4] ,
    \wbd_sdram_dat_i[3] ,
    \wbd_sdram_dat_i[2] ,
    \wbd_sdram_dat_i[1] ,
    \wbd_sdram_dat_i[0] }),
    .s1_wbd_dat_o({\wbd_sdram_dat_o[31] ,
    \wbd_sdram_dat_o[30] ,
    \wbd_sdram_dat_o[29] ,
    \wbd_sdram_dat_o[28] ,
    \wbd_sdram_dat_o[27] ,
    \wbd_sdram_dat_o[26] ,
    \wbd_sdram_dat_o[25] ,
    \wbd_sdram_dat_o[24] ,
    \wbd_sdram_dat_o[23] ,
    \wbd_sdram_dat_o[22] ,
    \wbd_sdram_dat_o[21] ,
    \wbd_sdram_dat_o[20] ,
    \wbd_sdram_dat_o[19] ,
    \wbd_sdram_dat_o[18] ,
    \wbd_sdram_dat_o[17] ,
    \wbd_sdram_dat_o[16] ,
    \wbd_sdram_dat_o[15] ,
    \wbd_sdram_dat_o[14] ,
    \wbd_sdram_dat_o[13] ,
    \wbd_sdram_dat_o[12] ,
    \wbd_sdram_dat_o[11] ,
    \wbd_sdram_dat_o[10] ,
    \wbd_sdram_dat_o[9] ,
    \wbd_sdram_dat_o[8] ,
    \wbd_sdram_dat_o[7] ,
    \wbd_sdram_dat_o[6] ,
    \wbd_sdram_dat_o[5] ,
    \wbd_sdram_dat_o[4] ,
    \wbd_sdram_dat_o[3] ,
    \wbd_sdram_dat_o[2] ,
    \wbd_sdram_dat_o[1] ,
    \wbd_sdram_dat_o[0] }),
    .s1_wbd_sel_o({\wbd_sdram_sel_o[3] ,
    \wbd_sdram_sel_o[2] ,
    \wbd_sdram_sel_o[1] ,
    \wbd_sdram_sel_o[0] }),
    .s2_wbd_adr_o({\wbd_glbl_adr_o[7] ,
    \wbd_glbl_adr_o[6] ,
    \wbd_glbl_adr_o[5] ,
    \wbd_glbl_adr_o[4] ,
    \wbd_glbl_adr_o[3] ,
    \wbd_glbl_adr_o[2] ,
    \wbd_glbl_adr_o[1] ,
    \wbd_glbl_adr_o[0] }),
    .s2_wbd_dat_i({\wbd_glbl_dat_i[31] ,
    \wbd_glbl_dat_i[30] ,
    \wbd_glbl_dat_i[29] ,
    \wbd_glbl_dat_i[28] ,
    \wbd_glbl_dat_i[27] ,
    \wbd_glbl_dat_i[26] ,
    \wbd_glbl_dat_i[25] ,
    \wbd_glbl_dat_i[24] ,
    \wbd_glbl_dat_i[23] ,
    \wbd_glbl_dat_i[22] ,
    \wbd_glbl_dat_i[21] ,
    \wbd_glbl_dat_i[20] ,
    \wbd_glbl_dat_i[19] ,
    \wbd_glbl_dat_i[18] ,
    \wbd_glbl_dat_i[17] ,
    \wbd_glbl_dat_i[16] ,
    \wbd_glbl_dat_i[15] ,
    \wbd_glbl_dat_i[14] ,
    \wbd_glbl_dat_i[13] ,
    \wbd_glbl_dat_i[12] ,
    \wbd_glbl_dat_i[11] ,
    \wbd_glbl_dat_i[10] ,
    \wbd_glbl_dat_i[9] ,
    \wbd_glbl_dat_i[8] ,
    \wbd_glbl_dat_i[7] ,
    \wbd_glbl_dat_i[6] ,
    \wbd_glbl_dat_i[5] ,
    \wbd_glbl_dat_i[4] ,
    \wbd_glbl_dat_i[3] ,
    \wbd_glbl_dat_i[2] ,
    \wbd_glbl_dat_i[1] ,
    \wbd_glbl_dat_i[0] }),
    .s2_wbd_dat_o({\wbd_glbl_dat_o[31] ,
    \wbd_glbl_dat_o[30] ,
    \wbd_glbl_dat_o[29] ,
    \wbd_glbl_dat_o[28] ,
    \wbd_glbl_dat_o[27] ,
    \wbd_glbl_dat_o[26] ,
    \wbd_glbl_dat_o[25] ,
    \wbd_glbl_dat_o[24] ,
    \wbd_glbl_dat_o[23] ,
    \wbd_glbl_dat_o[22] ,
    \wbd_glbl_dat_o[21] ,
    \wbd_glbl_dat_o[20] ,
    \wbd_glbl_dat_o[19] ,
    \wbd_glbl_dat_o[18] ,
    \wbd_glbl_dat_o[17] ,
    \wbd_glbl_dat_o[16] ,
    \wbd_glbl_dat_o[15] ,
    \wbd_glbl_dat_o[14] ,
    \wbd_glbl_dat_o[13] ,
    \wbd_glbl_dat_o[12] ,
    \wbd_glbl_dat_o[11] ,
    \wbd_glbl_dat_o[10] ,
    \wbd_glbl_dat_o[9] ,
    \wbd_glbl_dat_o[8] ,
    \wbd_glbl_dat_o[7] ,
    \wbd_glbl_dat_o[6] ,
    \wbd_glbl_dat_o[5] ,
    \wbd_glbl_dat_o[4] ,
    \wbd_glbl_dat_o[3] ,
    \wbd_glbl_dat_o[2] ,
    \wbd_glbl_dat_o[1] ,
    \wbd_glbl_dat_o[0] }),
    .s2_wbd_sel_o({\wbd_glbl_sel_o[3] ,
    \wbd_glbl_sel_o[2] ,
    \wbd_glbl_sel_o[1] ,
    \wbd_glbl_sel_o[0] }),
    .s3_wbd_adr_o({\wbd_uart_adr_o[7] ,
    \wbd_uart_adr_o[6] ,
    \wbd_uart_adr_o[5] ,
    \wbd_uart_adr_o[4] ,
    \wbd_uart_adr_o[3] ,
    \wbd_uart_adr_o[2] ,
    \wbd_uart_adr_o[1] ,
    \wbd_uart_adr_o[0] }),
    .s3_wbd_dat_i({\wbd_uart_dat_i[7] ,
    \wbd_uart_dat_i[6] ,
    \wbd_uart_dat_i[5] ,
    \wbd_uart_dat_i[4] ,
    \wbd_uart_dat_i[3] ,
    \wbd_uart_dat_i[2] ,
    \wbd_uart_dat_i[1] ,
    \wbd_uart_dat_i[0] }),
    .s3_wbd_dat_o({\wbd_uart_dat_o[7] ,
    \wbd_uart_dat_o[6] ,
    \wbd_uart_dat_o[5] ,
    \wbd_uart_dat_o[4] ,
    \wbd_uart_dat_o[3] ,
    \wbd_uart_dat_o[2] ,
    \wbd_uart_dat_o[1] ,
    \wbd_uart_dat_o[0] }));
 scr1_top_wb u_riscv_top (.core_clk(cpu_clk),
    .cpu_rst_n(cpu_rst_n),
    .pwrup_rst_n(wbd_int_rst_n),
    .rst_n(wbd_int_rst_n),
    .rtc_clk(rtc_clk),
    .soft_irq(soft_irq),
    .wb_clk(wbd_clk_riscv),
    .wb_rst_n(wbd_int_rst_n),
    .wbd_dmem_ack_i(wbd_riscv_dmem_ack_o),
    .wbd_dmem_err_i(wbd_riscv_dmem_err_o),
    .wbd_dmem_stb_o(wbd_riscv_dmem_stb_i),
    .wbd_dmem_we_o(wbd_riscv_dmem_we_i),
    .wbd_imem_ack_i(wbd_riscv_imem_ack_o),
    .wbd_imem_err_i(wbd_riscv_imem_err_o),
    .wbd_imem_stb_o(wbd_riscv_imem_stb_i),
    .wbd_imem_we_o(wbd_riscv_imem_we_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .fuse_mhartid({\fuse_mhartid[31] ,
    \fuse_mhartid[30] ,
    \fuse_mhartid[29] ,
    \fuse_mhartid[28] ,
    \fuse_mhartid[27] ,
    \fuse_mhartid[26] ,
    \fuse_mhartid[25] ,
    \fuse_mhartid[24] ,
    \fuse_mhartid[23] ,
    \fuse_mhartid[22] ,
    \fuse_mhartid[21] ,
    \fuse_mhartid[20] ,
    \fuse_mhartid[19] ,
    \fuse_mhartid[18] ,
    \fuse_mhartid[17] ,
    \fuse_mhartid[16] ,
    \fuse_mhartid[15] ,
    \fuse_mhartid[14] ,
    \fuse_mhartid[13] ,
    \fuse_mhartid[12] ,
    \fuse_mhartid[11] ,
    \fuse_mhartid[10] ,
    \fuse_mhartid[9] ,
    \fuse_mhartid[8] ,
    \fuse_mhartid[7] ,
    \fuse_mhartid[6] ,
    \fuse_mhartid[5] ,
    \fuse_mhartid[4] ,
    \fuse_mhartid[3] ,
    \fuse_mhartid[2] ,
    \fuse_mhartid[1] ,
    \fuse_mhartid[0] }),
    .irq_lines({\irq_lines[15] ,
    \irq_lines[14] ,
    \irq_lines[13] ,
    \irq_lines[12] ,
    \irq_lines[11] ,
    \irq_lines[10] ,
    \irq_lines[9] ,
    \irq_lines[8] ,
    \irq_lines[7] ,
    \irq_lines[6] ,
    \irq_lines[5] ,
    \irq_lines[4] ,
    \irq_lines[3] ,
    \irq_lines[2] ,
    \irq_lines[1] ,
    \irq_lines[0] }),
    .riscv_debug({la_data_out[63],
    la_data_out[62],
    la_data_out[61],
    la_data_out[60],
    la_data_out[59],
    la_data_out[58],
    la_data_out[57],
    la_data_out[56],
    la_data_out[55],
    la_data_out[54],
    la_data_out[53],
    la_data_out[52],
    la_data_out[51],
    la_data_out[50],
    la_data_out[49],
    la_data_out[48],
    la_data_out[47],
    la_data_out[46],
    la_data_out[45],
    la_data_out[44],
    la_data_out[43],
    la_data_out[42],
    la_data_out[41],
    la_data_out[40],
    la_data_out[39],
    la_data_out[38],
    la_data_out[37],
    la_data_out[36],
    la_data_out[35],
    la_data_out[34],
    la_data_out[33],
    la_data_out[32],
    la_data_out[31],
    la_data_out[30],
    la_data_out[29],
    la_data_out[28],
    la_data_out[27],
    la_data_out[26],
    la_data_out[25],
    la_data_out[24],
    la_data_out[23],
    la_data_out[22],
    la_data_out[21],
    la_data_out[20],
    la_data_out[19],
    la_data_out[18],
    la_data_out[17],
    la_data_out[16],
    la_data_out[15],
    la_data_out[14],
    la_data_out[13],
    la_data_out[12],
    la_data_out[11],
    la_data_out[10],
    la_data_out[9],
    la_data_out[8],
    la_data_out[7],
    la_data_out[6],
    la_data_out[5],
    la_data_out[4],
    la_data_out[3],
    la_data_out[2],
    la_data_out[1],
    la_data_out[0]}),
    .wbd_dmem_adr_o({\wbd_riscv_dmem_adr_i[31] ,
    \wbd_riscv_dmem_adr_i[30] ,
    \wbd_riscv_dmem_adr_i[29] ,
    \wbd_riscv_dmem_adr_i[28] ,
    \wbd_riscv_dmem_adr_i[27] ,
    \wbd_riscv_dmem_adr_i[26] ,
    \wbd_riscv_dmem_adr_i[25] ,
    \wbd_riscv_dmem_adr_i[24] ,
    \wbd_riscv_dmem_adr_i[23] ,
    \wbd_riscv_dmem_adr_i[22] ,
    \wbd_riscv_dmem_adr_i[21] ,
    \wbd_riscv_dmem_adr_i[20] ,
    \wbd_riscv_dmem_adr_i[19] ,
    \wbd_riscv_dmem_adr_i[18] ,
    \wbd_riscv_dmem_adr_i[17] ,
    \wbd_riscv_dmem_adr_i[16] ,
    \wbd_riscv_dmem_adr_i[15] ,
    \wbd_riscv_dmem_adr_i[14] ,
    \wbd_riscv_dmem_adr_i[13] ,
    \wbd_riscv_dmem_adr_i[12] ,
    \wbd_riscv_dmem_adr_i[11] ,
    \wbd_riscv_dmem_adr_i[10] ,
    \wbd_riscv_dmem_adr_i[9] ,
    \wbd_riscv_dmem_adr_i[8] ,
    \wbd_riscv_dmem_adr_i[7] ,
    \wbd_riscv_dmem_adr_i[6] ,
    \wbd_riscv_dmem_adr_i[5] ,
    \wbd_riscv_dmem_adr_i[4] ,
    \wbd_riscv_dmem_adr_i[3] ,
    \wbd_riscv_dmem_adr_i[2] ,
    \wbd_riscv_dmem_adr_i[1] ,
    \wbd_riscv_dmem_adr_i[0] }),
    .wbd_dmem_dat_i({\wbd_riscv_dmem_dat_o[31] ,
    \wbd_riscv_dmem_dat_o[30] ,
    \wbd_riscv_dmem_dat_o[29] ,
    \wbd_riscv_dmem_dat_o[28] ,
    \wbd_riscv_dmem_dat_o[27] ,
    \wbd_riscv_dmem_dat_o[26] ,
    \wbd_riscv_dmem_dat_o[25] ,
    \wbd_riscv_dmem_dat_o[24] ,
    \wbd_riscv_dmem_dat_o[23] ,
    \wbd_riscv_dmem_dat_o[22] ,
    \wbd_riscv_dmem_dat_o[21] ,
    \wbd_riscv_dmem_dat_o[20] ,
    \wbd_riscv_dmem_dat_o[19] ,
    \wbd_riscv_dmem_dat_o[18] ,
    \wbd_riscv_dmem_dat_o[17] ,
    \wbd_riscv_dmem_dat_o[16] ,
    \wbd_riscv_dmem_dat_o[15] ,
    \wbd_riscv_dmem_dat_o[14] ,
    \wbd_riscv_dmem_dat_o[13] ,
    \wbd_riscv_dmem_dat_o[12] ,
    \wbd_riscv_dmem_dat_o[11] ,
    \wbd_riscv_dmem_dat_o[10] ,
    \wbd_riscv_dmem_dat_o[9] ,
    \wbd_riscv_dmem_dat_o[8] ,
    \wbd_riscv_dmem_dat_o[7] ,
    \wbd_riscv_dmem_dat_o[6] ,
    \wbd_riscv_dmem_dat_o[5] ,
    \wbd_riscv_dmem_dat_o[4] ,
    \wbd_riscv_dmem_dat_o[3] ,
    \wbd_riscv_dmem_dat_o[2] ,
    \wbd_riscv_dmem_dat_o[1] ,
    \wbd_riscv_dmem_dat_o[0] }),
    .wbd_dmem_dat_o({\wbd_riscv_dmem_dat_i[31] ,
    \wbd_riscv_dmem_dat_i[30] ,
    \wbd_riscv_dmem_dat_i[29] ,
    \wbd_riscv_dmem_dat_i[28] ,
    \wbd_riscv_dmem_dat_i[27] ,
    \wbd_riscv_dmem_dat_i[26] ,
    \wbd_riscv_dmem_dat_i[25] ,
    \wbd_riscv_dmem_dat_i[24] ,
    \wbd_riscv_dmem_dat_i[23] ,
    \wbd_riscv_dmem_dat_i[22] ,
    \wbd_riscv_dmem_dat_i[21] ,
    \wbd_riscv_dmem_dat_i[20] ,
    \wbd_riscv_dmem_dat_i[19] ,
    \wbd_riscv_dmem_dat_i[18] ,
    \wbd_riscv_dmem_dat_i[17] ,
    \wbd_riscv_dmem_dat_i[16] ,
    \wbd_riscv_dmem_dat_i[15] ,
    \wbd_riscv_dmem_dat_i[14] ,
    \wbd_riscv_dmem_dat_i[13] ,
    \wbd_riscv_dmem_dat_i[12] ,
    \wbd_riscv_dmem_dat_i[11] ,
    \wbd_riscv_dmem_dat_i[10] ,
    \wbd_riscv_dmem_dat_i[9] ,
    \wbd_riscv_dmem_dat_i[8] ,
    \wbd_riscv_dmem_dat_i[7] ,
    \wbd_riscv_dmem_dat_i[6] ,
    \wbd_riscv_dmem_dat_i[5] ,
    \wbd_riscv_dmem_dat_i[4] ,
    \wbd_riscv_dmem_dat_i[3] ,
    \wbd_riscv_dmem_dat_i[2] ,
    \wbd_riscv_dmem_dat_i[1] ,
    \wbd_riscv_dmem_dat_i[0] }),
    .wbd_dmem_sel_o({\wbd_riscv_dmem_sel_i[3] ,
    \wbd_riscv_dmem_sel_i[2] ,
    \wbd_riscv_dmem_sel_i[1] ,
    \wbd_riscv_dmem_sel_i[0] }),
    .wbd_imem_adr_o({\wbd_riscv_imem_adr_i[31] ,
    \wbd_riscv_imem_adr_i[30] ,
    \wbd_riscv_imem_adr_i[29] ,
    \wbd_riscv_imem_adr_i[28] ,
    \wbd_riscv_imem_adr_i[27] ,
    \wbd_riscv_imem_adr_i[26] ,
    \wbd_riscv_imem_adr_i[25] ,
    \wbd_riscv_imem_adr_i[24] ,
    \wbd_riscv_imem_adr_i[23] ,
    \wbd_riscv_imem_adr_i[22] ,
    \wbd_riscv_imem_adr_i[21] ,
    \wbd_riscv_imem_adr_i[20] ,
    \wbd_riscv_imem_adr_i[19] ,
    \wbd_riscv_imem_adr_i[18] ,
    \wbd_riscv_imem_adr_i[17] ,
    \wbd_riscv_imem_adr_i[16] ,
    \wbd_riscv_imem_adr_i[15] ,
    \wbd_riscv_imem_adr_i[14] ,
    \wbd_riscv_imem_adr_i[13] ,
    \wbd_riscv_imem_adr_i[12] ,
    \wbd_riscv_imem_adr_i[11] ,
    \wbd_riscv_imem_adr_i[10] ,
    \wbd_riscv_imem_adr_i[9] ,
    \wbd_riscv_imem_adr_i[8] ,
    \wbd_riscv_imem_adr_i[7] ,
    \wbd_riscv_imem_adr_i[6] ,
    \wbd_riscv_imem_adr_i[5] ,
    \wbd_riscv_imem_adr_i[4] ,
    \wbd_riscv_imem_adr_i[3] ,
    \wbd_riscv_imem_adr_i[2] ,
    \wbd_riscv_imem_adr_i[1] ,
    \wbd_riscv_imem_adr_i[0] }),
    .wbd_imem_dat_i({\wbd_riscv_imem_dat_o[31] ,
    \wbd_riscv_imem_dat_o[30] ,
    \wbd_riscv_imem_dat_o[29] ,
    \wbd_riscv_imem_dat_o[28] ,
    \wbd_riscv_imem_dat_o[27] ,
    \wbd_riscv_imem_dat_o[26] ,
    \wbd_riscv_imem_dat_o[25] ,
    \wbd_riscv_imem_dat_o[24] ,
    \wbd_riscv_imem_dat_o[23] ,
    \wbd_riscv_imem_dat_o[22] ,
    \wbd_riscv_imem_dat_o[21] ,
    \wbd_riscv_imem_dat_o[20] ,
    \wbd_riscv_imem_dat_o[19] ,
    \wbd_riscv_imem_dat_o[18] ,
    \wbd_riscv_imem_dat_o[17] ,
    \wbd_riscv_imem_dat_o[16] ,
    \wbd_riscv_imem_dat_o[15] ,
    \wbd_riscv_imem_dat_o[14] ,
    \wbd_riscv_imem_dat_o[13] ,
    \wbd_riscv_imem_dat_o[12] ,
    \wbd_riscv_imem_dat_o[11] ,
    \wbd_riscv_imem_dat_o[10] ,
    \wbd_riscv_imem_dat_o[9] ,
    \wbd_riscv_imem_dat_o[8] ,
    \wbd_riscv_imem_dat_o[7] ,
    \wbd_riscv_imem_dat_o[6] ,
    \wbd_riscv_imem_dat_o[5] ,
    \wbd_riscv_imem_dat_o[4] ,
    \wbd_riscv_imem_dat_o[3] ,
    \wbd_riscv_imem_dat_o[2] ,
    \wbd_riscv_imem_dat_o[1] ,
    \wbd_riscv_imem_dat_o[0] }),
    .wbd_imem_dat_o({\wbd_riscv_imem_dat_i[31] ,
    \wbd_riscv_imem_dat_i[30] ,
    \wbd_riscv_imem_dat_i[29] ,
    \wbd_riscv_imem_dat_i[28] ,
    \wbd_riscv_imem_dat_i[27] ,
    \wbd_riscv_imem_dat_i[26] ,
    \wbd_riscv_imem_dat_i[25] ,
    \wbd_riscv_imem_dat_i[24] ,
    \wbd_riscv_imem_dat_i[23] ,
    \wbd_riscv_imem_dat_i[22] ,
    \wbd_riscv_imem_dat_i[21] ,
    \wbd_riscv_imem_dat_i[20] ,
    \wbd_riscv_imem_dat_i[19] ,
    \wbd_riscv_imem_dat_i[18] ,
    \wbd_riscv_imem_dat_i[17] ,
    \wbd_riscv_imem_dat_i[16] ,
    \wbd_riscv_imem_dat_i[15] ,
    \wbd_riscv_imem_dat_i[14] ,
    \wbd_riscv_imem_dat_i[13] ,
    \wbd_riscv_imem_dat_i[12] ,
    \wbd_riscv_imem_dat_i[11] ,
    \wbd_riscv_imem_dat_i[10] ,
    \wbd_riscv_imem_dat_i[9] ,
    \wbd_riscv_imem_dat_i[8] ,
    \wbd_riscv_imem_dat_i[7] ,
    \wbd_riscv_imem_dat_i[6] ,
    \wbd_riscv_imem_dat_i[5] ,
    \wbd_riscv_imem_dat_i[4] ,
    \wbd_riscv_imem_dat_i[3] ,
    \wbd_riscv_imem_dat_i[2] ,
    \wbd_riscv_imem_dat_i[1] ,
    \wbd_riscv_imem_dat_i[0] }),
    .wbd_imem_sel_o({\wbd_riscv_imem_sel_i[3] ,
    \wbd_riscv_imem_sel_i[2] ,
    \wbd_riscv_imem_sel_i[1] ,
    \wbd_riscv_imem_sel_i[0] }));
 sdrc_top u_sdram_ctrl (.cfg_sdr_en(cfg_sdr_en),
    .sdr_init_done(sdr_init_done),
    .sdram_clk(sdram_clk),
    .sdram_resetn(sdram_rst_n),
    .wb_ack_o(wbd_sdram_ack_i),
    .wb_clk_i(wbd_clk_sdram),
    .wb_cyc_i(wbd_sdram_cyc_o),
    .wb_rst_n(wbd_int_rst_n),
    .wb_stb_i(wbd_sdram_stb_o),
    .wb_we_i(wbd_sdram_we_o),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .cfg_colbits({\cfg_colbits[1] ,
    \cfg_colbits[0] }),
    .cfg_req_depth({\cfg_req_depth[1] ,
    \cfg_req_depth[0] }),
    .cfg_sdr_cas({\cfg_sdr_cas[2] ,
    \cfg_sdr_cas[1] ,
    \cfg_sdr_cas[0] }),
    .cfg_sdr_mode_reg({\cfg_sdr_mode_reg[12] ,
    \cfg_sdr_mode_reg[11] ,
    \cfg_sdr_mode_reg[10] ,
    \cfg_sdr_mode_reg[9] ,
    \cfg_sdr_mode_reg[8] ,
    \cfg_sdr_mode_reg[7] ,
    \cfg_sdr_mode_reg[6] ,
    \cfg_sdr_mode_reg[5] ,
    \cfg_sdr_mode_reg[4] ,
    \cfg_sdr_mode_reg[3] ,
    \cfg_sdr_mode_reg[2] ,
    \cfg_sdr_mode_reg[1] ,
    \cfg_sdr_mode_reg[0] }),
    .cfg_sdr_rfmax({\cfg_sdr_rfmax[2] ,
    \cfg_sdr_rfmax[1] ,
    \cfg_sdr_rfmax[0] }),
    .cfg_sdr_rfsh({\cfg_sdr_rfsh[11] ,
    \cfg_sdr_rfsh[10] ,
    \cfg_sdr_rfsh[9] ,
    \cfg_sdr_rfsh[8] ,
    \cfg_sdr_rfsh[7] ,
    \cfg_sdr_rfsh[6] ,
    \cfg_sdr_rfsh[5] ,
    \cfg_sdr_rfsh[4] ,
    \cfg_sdr_rfsh[3] ,
    \cfg_sdr_rfsh[2] ,
    \cfg_sdr_rfsh[1] ,
    \cfg_sdr_rfsh[0] }),
    .cfg_sdr_tras_d({\cfg_sdr_tras_d[3] ,
    \cfg_sdr_tras_d[2] ,
    \cfg_sdr_tras_d[1] ,
    \cfg_sdr_tras_d[0] }),
    .cfg_sdr_trcar_d({\cfg_sdr_trcar_d[3] ,
    \cfg_sdr_trcar_d[2] ,
    \cfg_sdr_trcar_d[1] ,
    \cfg_sdr_trcar_d[0] }),
    .cfg_sdr_trcd_d({\cfg_sdr_trcd_d[3] ,
    \cfg_sdr_trcd_d[2] ,
    \cfg_sdr_trcd_d[1] ,
    \cfg_sdr_trcd_d[0] }),
    .cfg_sdr_trp_d({\cfg_sdr_trp_d[3] ,
    \cfg_sdr_trp_d[2] ,
    \cfg_sdr_trp_d[1] ,
    \cfg_sdr_trp_d[0] }),
    .cfg_sdr_twr_d({\cfg_sdr_twr_d[3] ,
    \cfg_sdr_twr_d[2] ,
    \cfg_sdr_twr_d[1] ,
    \cfg_sdr_twr_d[0] }),
    .cfg_sdr_width({\cfg_sdr_width[1] ,
    \cfg_sdr_width[0] }),
    .io_in({io_in_29_,
    io_in[28],
    io_in[27],
    io_in[26],
    io_in[25],
    io_in[24],
    io_in[23],
    io_in[22],
    io_in[21],
    io_in[20],
    io_in[19],
    io_in[18],
    io_in[17],
    io_in[16],
    io_in[15],
    io_in[14],
    io_in[13],
    io_in[12],
    io_in[11],
    io_in[10],
    io_in[9],
    io_in[8],
    io_in[7],
    io_in[6],
    io_in[5],
    io_in[4],
    io_in[3],
    io_in[2],
    io_in[1],
    io_in[0]}),
    .io_oeb({io_oeb[29],
    io_oeb[28],
    io_oeb[27],
    io_oeb[26],
    io_oeb[25],
    io_oeb[24],
    io_oeb[23],
    io_oeb[22],
    io_oeb[21],
    io_oeb[20],
    io_oeb[19],
    io_oeb[18],
    io_oeb[17],
    io_oeb[16],
    io_oeb[15],
    io_oeb[14],
    io_oeb[13],
    io_oeb[12],
    io_oeb[11],
    io_oeb[10],
    io_oeb[9],
    io_oeb[8],
    io_oeb[7],
    io_oeb[6],
    io_oeb[5],
    io_oeb[4],
    io_oeb[3],
    io_oeb[2],
    io_oeb[1],
    io_oeb[0]}),
    .io_out({io_out_29_,
    io_out[28],
    io_out[27],
    io_out[26],
    io_out[25],
    io_out[24],
    io_out[23],
    io_out[22],
    io_out[21],
    io_out[20],
    io_out[19],
    io_out[18],
    io_out[17],
    io_out[16],
    io_out[15],
    io_out[14],
    io_out[13],
    io_out[12],
    io_out[11],
    io_out[10],
    io_out[9],
    io_out[8],
    io_out[7],
    io_out[6],
    io_out[5],
    io_out[4],
    io_out[3],
    io_out[2],
    io_out[1],
    io_out[0]}),
    .sdram_debug({la_data_out[127],
    la_data_out[126],
    la_data_out[125],
    la_data_out[124],
    la_data_out[123],
    la_data_out[122],
    la_data_out[121],
    la_data_out[120],
    la_data_out[119],
    la_data_out[118],
    la_data_out[117],
    la_data_out[116],
    la_data_out[115],
    la_data_out[114],
    la_data_out[113],
    la_data_out[112],
    la_data_out[111],
    la_data_out[110],
    la_data_out[109],
    la_data_out[108],
    la_data_out[107],
    la_data_out[106],
    la_data_out[105],
    la_data_out[104],
    la_data_out[103],
    la_data_out[102],
    la_data_out[101],
    la_data_out[100],
    la_data_out[99],
    la_data_out[98],
    la_data_out[97],
    la_data_out[96]}),
    .wb_addr_i({\wbd_sdram_adr_o[31] ,
    \wbd_sdram_adr_o[30] ,
    \wbd_sdram_adr_o[29] ,
    \wbd_sdram_adr_o[28] ,
    \wbd_sdram_adr_o[27] ,
    \wbd_sdram_adr_o[26] ,
    \wbd_sdram_adr_o[25] ,
    \wbd_sdram_adr_o[24] ,
    \wbd_sdram_adr_o[23] ,
    \wbd_sdram_adr_o[22] ,
    \wbd_sdram_adr_o[21] ,
    \wbd_sdram_adr_o[20] ,
    \wbd_sdram_adr_o[19] ,
    \wbd_sdram_adr_o[18] ,
    \wbd_sdram_adr_o[17] ,
    \wbd_sdram_adr_o[16] ,
    \wbd_sdram_adr_o[15] ,
    \wbd_sdram_adr_o[14] ,
    \wbd_sdram_adr_o[13] ,
    \wbd_sdram_adr_o[12] ,
    \wbd_sdram_adr_o[11] ,
    \wbd_sdram_adr_o[10] ,
    \wbd_sdram_adr_o[9] ,
    \wbd_sdram_adr_o[8] ,
    \wbd_sdram_adr_o[7] ,
    \wbd_sdram_adr_o[6] ,
    \wbd_sdram_adr_o[5] ,
    \wbd_sdram_adr_o[4] ,
    \wbd_sdram_adr_o[3] ,
    \wbd_sdram_adr_o[2] ,
    \wbd_sdram_adr_o[1] ,
    \wbd_sdram_adr_o[0] }),
    .wb_dat_i({\wbd_sdram_dat_o[31] ,
    \wbd_sdram_dat_o[30] ,
    \wbd_sdram_dat_o[29] ,
    \wbd_sdram_dat_o[28] ,
    \wbd_sdram_dat_o[27] ,
    \wbd_sdram_dat_o[26] ,
    \wbd_sdram_dat_o[25] ,
    \wbd_sdram_dat_o[24] ,
    \wbd_sdram_dat_o[23] ,
    \wbd_sdram_dat_o[22] ,
    \wbd_sdram_dat_o[21] ,
    \wbd_sdram_dat_o[20] ,
    \wbd_sdram_dat_o[19] ,
    \wbd_sdram_dat_o[18] ,
    \wbd_sdram_dat_o[17] ,
    \wbd_sdram_dat_o[16] ,
    \wbd_sdram_dat_o[15] ,
    \wbd_sdram_dat_o[14] ,
    \wbd_sdram_dat_o[13] ,
    \wbd_sdram_dat_o[12] ,
    \wbd_sdram_dat_o[11] ,
    \wbd_sdram_dat_o[10] ,
    \wbd_sdram_dat_o[9] ,
    \wbd_sdram_dat_o[8] ,
    \wbd_sdram_dat_o[7] ,
    \wbd_sdram_dat_o[6] ,
    \wbd_sdram_dat_o[5] ,
    \wbd_sdram_dat_o[4] ,
    \wbd_sdram_dat_o[3] ,
    \wbd_sdram_dat_o[2] ,
    \wbd_sdram_dat_o[1] ,
    \wbd_sdram_dat_o[0] }),
    .wb_dat_o({\wbd_sdram_dat_i[31] ,
    \wbd_sdram_dat_i[30] ,
    \wbd_sdram_dat_i[29] ,
    \wbd_sdram_dat_i[28] ,
    \wbd_sdram_dat_i[27] ,
    \wbd_sdram_dat_i[26] ,
    \wbd_sdram_dat_i[25] ,
    \wbd_sdram_dat_i[24] ,
    \wbd_sdram_dat_i[23] ,
    \wbd_sdram_dat_i[22] ,
    \wbd_sdram_dat_i[21] ,
    \wbd_sdram_dat_i[20] ,
    \wbd_sdram_dat_i[19] ,
    \wbd_sdram_dat_i[18] ,
    \wbd_sdram_dat_i[17] ,
    \wbd_sdram_dat_i[16] ,
    \wbd_sdram_dat_i[15] ,
    \wbd_sdram_dat_i[14] ,
    \wbd_sdram_dat_i[13] ,
    \wbd_sdram_dat_i[12] ,
    \wbd_sdram_dat_i[11] ,
    \wbd_sdram_dat_i[10] ,
    \wbd_sdram_dat_i[9] ,
    \wbd_sdram_dat_i[8] ,
    \wbd_sdram_dat_i[7] ,
    \wbd_sdram_dat_i[6] ,
    \wbd_sdram_dat_i[5] ,
    \wbd_sdram_dat_i[4] ,
    \wbd_sdram_dat_i[3] ,
    \wbd_sdram_dat_i[2] ,
    \wbd_sdram_dat_i[1] ,
    \wbd_sdram_dat_i[0] }),
    .wb_sel_i({\wbd_sdram_sel_o[3] ,
    \wbd_sdram_sel_o[2] ,
    \wbd_sdram_sel_o[1] ,
    \wbd_sdram_sel_o[0] }));
 clk_skew_adjust u_skew_glbl (.clk_in(wbd_clk_int),
    .clk_out(wbd_clk_glbl),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .sel({\cfg_clk_ctrl1[23] ,
    \cfg_clk_ctrl1[22] ,
    \cfg_clk_ctrl1[21] ,
    \cfg_clk_ctrl1[20] }));
 clk_skew_adjust u_skew_riscv (.clk_in(wbd_clk_int),
    .clk_out(wbd_clk_riscv),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .sel({\cfg_clk_ctrl1[7] ,
    \cfg_clk_ctrl1[6] ,
    \cfg_clk_ctrl1[5] ,
    \cfg_clk_ctrl1[4] }));
 clk_skew_adjust u_skew_sd_ci (.clk_in(io_in[29]),
    .clk_out(io_in_29_),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .sel({\cfg_clk_ctrl2[7] ,
    \cfg_clk_ctrl2[6] ,
    \cfg_clk_ctrl2[5] ,
    \cfg_clk_ctrl2[4] }));
 clk_skew_adjust u_skew_sd_co (.clk_in(sdram_clk),
    .clk_out(io_out[29]),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .sel({\cfg_clk_ctrl2[3] ,
    \cfg_clk_ctrl2[2] ,
    \cfg_clk_ctrl2[1] ,
    \cfg_clk_ctrl2[0] }));
 clk_skew_adjust u_skew_sdram (.clk_in(wbd_clk_int),
    .clk_out(wbd_clk_sdram),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .sel({\cfg_clk_ctrl1[19] ,
    \cfg_clk_ctrl1[18] ,
    \cfg_clk_ctrl1[17] ,
    \cfg_clk_ctrl1[16] }));
 clk_skew_adjust u_skew_sp_co (.clk_in(io_in_30_),
    .clk_out(io_out[30]),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .sel({\cfg_clk_ctrl2[11] ,
    \cfg_clk_ctrl2[10] ,
    \cfg_clk_ctrl2[9] ,
    \cfg_clk_ctrl2[8] }));
 clk_skew_adjust u_skew_spi (.clk_in(wbd_clk_int),
    .clk_out(wbd_clk_spi),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .sel({\cfg_clk_ctrl1[15] ,
    \cfg_clk_ctrl1[14] ,
    \cfg_clk_ctrl1[13] ,
    \cfg_clk_ctrl1[12] }));
 clk_skew_adjust u_skew_uart (.clk_in(wbd_clk_int),
    .clk_out(wbd_clk_uart),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .sel({\cfg_clk_ctrl1[11] ,
    \cfg_clk_ctrl1[10] ,
    \cfg_clk_ctrl1[9] ,
    \cfg_clk_ctrl1[8] }));
 clk_skew_adjust u_skew_wh (.clk_in(wbd_clk_int),
    .clk_out(wbd_clk_wh),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .sel({\cfg_clk_ctrl1[27] ,
    \cfg_clk_ctrl1[26] ,
    \cfg_clk_ctrl1[25] ,
    \cfg_clk_ctrl1[24] }));
 clk_skew_adjust u_skew_wi (.clk_in(wbd_clk_int),
    .clk_out(wbd_clk_wi),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .sel({\cfg_clk_ctrl1[3] ,
    \cfg_clk_ctrl1[2] ,
    \cfg_clk_ctrl1[1] ,
    \cfg_clk_ctrl1[0] }));
 spim_top u_spi_master (.mclk(wbd_clk_spi),
    .rst_n(spi_rst_n),
    .wbd_ack_o(wbd_spim_ack_i),
    .wbd_err_o(wbd_spim_err_i),
    .wbd_stb_i(wbd_spim_stb_o),
    .wbd_we_i(wbd_spim_we_o),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({io_in[35],
    io_in[34],
    io_in[33],
    io_in[32]}),
    .io_oeb({io_oeb[35],
    io_oeb[34],
    io_oeb[33],
    io_oeb[32],
    io_oeb[31],
    io_oeb[30]}),
    .io_out({io_out[35],
    io_out[34],
    io_out[33],
    io_out[32],
    io_out[31],
    io_in_30_}),
    .spi_debug({la_data_out[95],
    la_data_out[94],
    la_data_out[93],
    la_data_out[92],
    la_data_out[91],
    la_data_out[90],
    la_data_out[89],
    la_data_out[88],
    la_data_out[87],
    la_data_out[86],
    la_data_out[85],
    la_data_out[84],
    la_data_out[83],
    la_data_out[82],
    la_data_out[81],
    la_data_out[80],
    la_data_out[79],
    la_data_out[78],
    la_data_out[77],
    la_data_out[76],
    la_data_out[75],
    la_data_out[74],
    la_data_out[73],
    la_data_out[72],
    la_data_out[71],
    la_data_out[70],
    la_data_out[69],
    la_data_out[68],
    la_data_out[67],
    la_data_out[66],
    la_data_out[65],
    la_data_out[64]}),
    .wbd_adr_i({\wbd_spim_adr_o[31] ,
    \wbd_spim_adr_o[30] ,
    \wbd_spim_adr_o[29] ,
    \wbd_spim_adr_o[28] ,
    \wbd_spim_adr_o[27] ,
    \wbd_spim_adr_o[26] ,
    \wbd_spim_adr_o[25] ,
    \wbd_spim_adr_o[24] ,
    \wbd_spim_adr_o[23] ,
    \wbd_spim_adr_o[22] ,
    \wbd_spim_adr_o[21] ,
    \wbd_spim_adr_o[20] ,
    \wbd_spim_adr_o[19] ,
    \wbd_spim_adr_o[18] ,
    \wbd_spim_adr_o[17] ,
    \wbd_spim_adr_o[16] ,
    \wbd_spim_adr_o[15] ,
    \wbd_spim_adr_o[14] ,
    \wbd_spim_adr_o[13] ,
    \wbd_spim_adr_o[12] ,
    \wbd_spim_adr_o[11] ,
    \wbd_spim_adr_o[10] ,
    \wbd_spim_adr_o[9] ,
    \wbd_spim_adr_o[8] ,
    \wbd_spim_adr_o[7] ,
    \wbd_spim_adr_o[6] ,
    \wbd_spim_adr_o[5] ,
    \wbd_spim_adr_o[4] ,
    \wbd_spim_adr_o[3] ,
    \wbd_spim_adr_o[2] ,
    \wbd_spim_adr_o[1] ,
    \wbd_spim_adr_o[0] }),
    .wbd_dat_i({\wbd_spim_dat_o[31] ,
    \wbd_spim_dat_o[30] ,
    \wbd_spim_dat_o[29] ,
    \wbd_spim_dat_o[28] ,
    \wbd_spim_dat_o[27] ,
    \wbd_spim_dat_o[26] ,
    \wbd_spim_dat_o[25] ,
    \wbd_spim_dat_o[24] ,
    \wbd_spim_dat_o[23] ,
    \wbd_spim_dat_o[22] ,
    \wbd_spim_dat_o[21] ,
    \wbd_spim_dat_o[20] ,
    \wbd_spim_dat_o[19] ,
    \wbd_spim_dat_o[18] ,
    \wbd_spim_dat_o[17] ,
    \wbd_spim_dat_o[16] ,
    \wbd_spim_dat_o[15] ,
    \wbd_spim_dat_o[14] ,
    \wbd_spim_dat_o[13] ,
    \wbd_spim_dat_o[12] ,
    \wbd_spim_dat_o[11] ,
    \wbd_spim_dat_o[10] ,
    \wbd_spim_dat_o[9] ,
    \wbd_spim_dat_o[8] ,
    \wbd_spim_dat_o[7] ,
    \wbd_spim_dat_o[6] ,
    \wbd_spim_dat_o[5] ,
    \wbd_spim_dat_o[4] ,
    \wbd_spim_dat_o[3] ,
    \wbd_spim_dat_o[2] ,
    \wbd_spim_dat_o[1] ,
    \wbd_spim_dat_o[0] }),
    .wbd_dat_o({\wbd_spim_dat_i[31] ,
    \wbd_spim_dat_i[30] ,
    \wbd_spim_dat_i[29] ,
    \wbd_spim_dat_i[28] ,
    \wbd_spim_dat_i[27] ,
    \wbd_spim_dat_i[26] ,
    \wbd_spim_dat_i[25] ,
    \wbd_spim_dat_i[24] ,
    \wbd_spim_dat_i[23] ,
    \wbd_spim_dat_i[22] ,
    \wbd_spim_dat_i[21] ,
    \wbd_spim_dat_i[20] ,
    \wbd_spim_dat_i[19] ,
    \wbd_spim_dat_i[18] ,
    \wbd_spim_dat_i[17] ,
    \wbd_spim_dat_i[16] ,
    \wbd_spim_dat_i[15] ,
    \wbd_spim_dat_i[14] ,
    \wbd_spim_dat_i[13] ,
    \wbd_spim_dat_i[12] ,
    \wbd_spim_dat_i[11] ,
    \wbd_spim_dat_i[10] ,
    \wbd_spim_dat_i[9] ,
    \wbd_spim_dat_i[8] ,
    \wbd_spim_dat_i[7] ,
    \wbd_spim_dat_i[6] ,
    \wbd_spim_dat_i[5] ,
    \wbd_spim_dat_i[4] ,
    \wbd_spim_dat_i[3] ,
    \wbd_spim_dat_i[2] ,
    \wbd_spim_dat_i[1] ,
    \wbd_spim_dat_i[0] }),
    .wbd_sel_i({\wbd_spim_sel_o[3] ,
    \wbd_spim_sel_o[2] ,
    \wbd_spim_sel_o[1] ,
    \wbd_spim_sel_o[0] }));
 uart_core u_uart_core (.app_clk(wbd_clk_uart),
    .arst_n(wbd_int_rst_n),
    .reg_ack(wbd_uart_ack_i),
    .reg_be(wbd_uart_sel_o),
    .reg_cs(wbd_uart_stb_o),
    .reg_wr(wbd_uart_we_o),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({io_in[37],
    io_in[36]}),
    .io_oeb({io_oeb[37],
    io_oeb[36]}),
    .io_out({io_out[37],
    io_out[36]}),
    .reg_addr({\wbd_uart_adr_o[5] ,
    \wbd_uart_adr_o[4] ,
    \wbd_uart_adr_o[3] ,
    \wbd_uart_adr_o[2] }),
    .reg_rdata({\wbd_uart_dat_i[7] ,
    \wbd_uart_dat_i[6] ,
    \wbd_uart_dat_i[5] ,
    \wbd_uart_dat_i[4] ,
    \wbd_uart_dat_i[3] ,
    \wbd_uart_dat_i[2] ,
    \wbd_uart_dat_i[1] ,
    \wbd_uart_dat_i[0] }),
    .reg_wdata({\wbd_uart_dat_o[7] ,
    \wbd_uart_dat_o[6] ,
    \wbd_uart_dat_o[5] ,
    \wbd_uart_dat_o[4] ,
    \wbd_uart_dat_o[3] ,
    \wbd_uart_dat_o[2] ,
    \wbd_uart_dat_o[1] ,
    \wbd_uart_dat_o[0] }));
 wb_host u_wb_host (.cpu_clk(cpu_clk),
    .cpu_rst_n(cpu_rst_n),
    .rtc_clk(rtc_clk),
    .sdram_clk(sdram_clk),
    .sdram_rst_n(sdram_rst_n),
    .spi_rst_n(spi_rst_n),
    .user_clock1(wb_clk_i),
    .user_clock2(user_clock2),
    .wbd_int_rst_n(wbd_int_rst_n),
    .wbm_ack_o(wbs_ack_o),
    .wbm_clk_i(wb_clk_i),
    .wbm_cyc_i(wbs_cyc_i),
    .wbm_rst_i(wb_rst_i),
    .wbm_stb_i(wbs_stb_i),
    .wbm_we_i(wbs_we_i),
    .wbs_ack_i(wbd_int_ack_o),
    .wbs_clk_i(wbd_clk_wh),
    .wbs_clk_out(wbd_clk_int),
    .wbs_cyc_o(wbd_int_cyc_i),
    .wbs_err_i(wbd_int_err_o),
    .wbs_stb_o(wbd_int_stb_i),
    .wbs_we_o(wbd_int_we_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .cfg_clk_ctrl1({\cfg_clk_ctrl1[31] ,
    \cfg_clk_ctrl1[30] ,
    \cfg_clk_ctrl1[29] ,
    \cfg_clk_ctrl1[28] ,
    \cfg_clk_ctrl1[27] ,
    \cfg_clk_ctrl1[26] ,
    \cfg_clk_ctrl1[25] ,
    \cfg_clk_ctrl1[24] ,
    \cfg_clk_ctrl1[23] ,
    \cfg_clk_ctrl1[22] ,
    \cfg_clk_ctrl1[21] ,
    \cfg_clk_ctrl1[20] ,
    \cfg_clk_ctrl1[19] ,
    \cfg_clk_ctrl1[18] ,
    \cfg_clk_ctrl1[17] ,
    \cfg_clk_ctrl1[16] ,
    \cfg_clk_ctrl1[15] ,
    \cfg_clk_ctrl1[14] ,
    \cfg_clk_ctrl1[13] ,
    \cfg_clk_ctrl1[12] ,
    \cfg_clk_ctrl1[11] ,
    \cfg_clk_ctrl1[10] ,
    \cfg_clk_ctrl1[9] ,
    \cfg_clk_ctrl1[8] ,
    \cfg_clk_ctrl1[7] ,
    \cfg_clk_ctrl1[6] ,
    \cfg_clk_ctrl1[5] ,
    \cfg_clk_ctrl1[4] ,
    \cfg_clk_ctrl1[3] ,
    \cfg_clk_ctrl1[2] ,
    \cfg_clk_ctrl1[1] ,
    \cfg_clk_ctrl1[0] }),
    .cfg_clk_ctrl2({\cfg_clk_ctrl2[31] ,
    \cfg_clk_ctrl2[30] ,
    \cfg_clk_ctrl2[29] ,
    \cfg_clk_ctrl2[28] ,
    \cfg_clk_ctrl2[27] ,
    \cfg_clk_ctrl2[26] ,
    \cfg_clk_ctrl2[25] ,
    \cfg_clk_ctrl2[24] ,
    \cfg_clk_ctrl2[23] ,
    \cfg_clk_ctrl2[22] ,
    \cfg_clk_ctrl2[21] ,
    \cfg_clk_ctrl2[20] ,
    \cfg_clk_ctrl2[19] ,
    \cfg_clk_ctrl2[18] ,
    \cfg_clk_ctrl2[17] ,
    \cfg_clk_ctrl2[16] ,
    \cfg_clk_ctrl2[15] ,
    \cfg_clk_ctrl2[14] ,
    \cfg_clk_ctrl2[13] ,
    \cfg_clk_ctrl2[12] ,
    \cfg_clk_ctrl2[11] ,
    \cfg_clk_ctrl2[10] ,
    \cfg_clk_ctrl2[9] ,
    \cfg_clk_ctrl2[8] ,
    \cfg_clk_ctrl2[7] ,
    \cfg_clk_ctrl2[6] ,
    \cfg_clk_ctrl2[5] ,
    \cfg_clk_ctrl2[4] ,
    \cfg_clk_ctrl2[3] ,
    \cfg_clk_ctrl2[2] ,
    \cfg_clk_ctrl2[1] ,
    \cfg_clk_ctrl2[0] }),
    .wbm_adr_i({wbs_adr_i[31],
    wbs_adr_i[30],
    wbs_adr_i[29],
    wbs_adr_i[28],
    wbs_adr_i[27],
    wbs_adr_i[26],
    wbs_adr_i[25],
    wbs_adr_i[24],
    wbs_adr_i[23],
    wbs_adr_i[22],
    wbs_adr_i[21],
    wbs_adr_i[20],
    wbs_adr_i[19],
    wbs_adr_i[18],
    wbs_adr_i[17],
    wbs_adr_i[16],
    wbs_adr_i[15],
    wbs_adr_i[14],
    wbs_adr_i[13],
    wbs_adr_i[12],
    wbs_adr_i[11],
    wbs_adr_i[10],
    wbs_adr_i[9],
    wbs_adr_i[8],
    wbs_adr_i[7],
    wbs_adr_i[6],
    wbs_adr_i[5],
    wbs_adr_i[4],
    wbs_adr_i[3],
    wbs_adr_i[2],
    wbs_adr_i[1],
    wbs_adr_i[0]}),
    .wbm_dat_i({wbs_dat_i[31],
    wbs_dat_i[30],
    wbs_dat_i[29],
    wbs_dat_i[28],
    wbs_dat_i[27],
    wbs_dat_i[26],
    wbs_dat_i[25],
    wbs_dat_i[24],
    wbs_dat_i[23],
    wbs_dat_i[22],
    wbs_dat_i[21],
    wbs_dat_i[20],
    wbs_dat_i[19],
    wbs_dat_i[18],
    wbs_dat_i[17],
    wbs_dat_i[16],
    wbs_dat_i[15],
    wbs_dat_i[14],
    wbs_dat_i[13],
    wbs_dat_i[12],
    wbs_dat_i[11],
    wbs_dat_i[10],
    wbs_dat_i[9],
    wbs_dat_i[8],
    wbs_dat_i[7],
    wbs_dat_i[6],
    wbs_dat_i[5],
    wbs_dat_i[4],
    wbs_dat_i[3],
    wbs_dat_i[2],
    wbs_dat_i[1],
    wbs_dat_i[0]}),
    .wbm_dat_o({wbs_dat_o[31],
    wbs_dat_o[30],
    wbs_dat_o[29],
    wbs_dat_o[28],
    wbs_dat_o[27],
    wbs_dat_o[26],
    wbs_dat_o[25],
    wbs_dat_o[24],
    wbs_dat_o[23],
    wbs_dat_o[22],
    wbs_dat_o[21],
    wbs_dat_o[20],
    wbs_dat_o[19],
    wbs_dat_o[18],
    wbs_dat_o[17],
    wbs_dat_o[16],
    wbs_dat_o[15],
    wbs_dat_o[14],
    wbs_dat_o[13],
    wbs_dat_o[12],
    wbs_dat_o[11],
    wbs_dat_o[10],
    wbs_dat_o[9],
    wbs_dat_o[8],
    wbs_dat_o[7],
    wbs_dat_o[6],
    wbs_dat_o[5],
    wbs_dat_o[4],
    wbs_dat_o[3],
    wbs_dat_o[2],
    wbs_dat_o[1],
    wbs_dat_o[0]}),
    .wbm_sel_i({wbs_sel_i[3],
    wbs_sel_i[2],
    wbs_sel_i[1],
    wbs_sel_i[0]}),
    .wbs_adr_o({\wbd_int_adr_i[31] ,
    \wbd_int_adr_i[30] ,
    \wbd_int_adr_i[29] ,
    \wbd_int_adr_i[28] ,
    \wbd_int_adr_i[27] ,
    \wbd_int_adr_i[26] ,
    \wbd_int_adr_i[25] ,
    \wbd_int_adr_i[24] ,
    \wbd_int_adr_i[23] ,
    \wbd_int_adr_i[22] ,
    \wbd_int_adr_i[21] ,
    \wbd_int_adr_i[20] ,
    \wbd_int_adr_i[19] ,
    \wbd_int_adr_i[18] ,
    \wbd_int_adr_i[17] ,
    \wbd_int_adr_i[16] ,
    \wbd_int_adr_i[15] ,
    \wbd_int_adr_i[14] ,
    \wbd_int_adr_i[13] ,
    \wbd_int_adr_i[12] ,
    \wbd_int_adr_i[11] ,
    \wbd_int_adr_i[10] ,
    \wbd_int_adr_i[9] ,
    \wbd_int_adr_i[8] ,
    \wbd_int_adr_i[7] ,
    \wbd_int_adr_i[6] ,
    \wbd_int_adr_i[5] ,
    \wbd_int_adr_i[4] ,
    \wbd_int_adr_i[3] ,
    \wbd_int_adr_i[2] ,
    \wbd_int_adr_i[1] ,
    \wbd_int_adr_i[0] }),
    .wbs_dat_i({\wbd_int_dat_o[31] ,
    \wbd_int_dat_o[30] ,
    \wbd_int_dat_o[29] ,
    \wbd_int_dat_o[28] ,
    \wbd_int_dat_o[27] ,
    \wbd_int_dat_o[26] ,
    \wbd_int_dat_o[25] ,
    \wbd_int_dat_o[24] ,
    \wbd_int_dat_o[23] ,
    \wbd_int_dat_o[22] ,
    \wbd_int_dat_o[21] ,
    \wbd_int_dat_o[20] ,
    \wbd_int_dat_o[19] ,
    \wbd_int_dat_o[18] ,
    \wbd_int_dat_o[17] ,
    \wbd_int_dat_o[16] ,
    \wbd_int_dat_o[15] ,
    \wbd_int_dat_o[14] ,
    \wbd_int_dat_o[13] ,
    \wbd_int_dat_o[12] ,
    \wbd_int_dat_o[11] ,
    \wbd_int_dat_o[10] ,
    \wbd_int_dat_o[9] ,
    \wbd_int_dat_o[8] ,
    \wbd_int_dat_o[7] ,
    \wbd_int_dat_o[6] ,
    \wbd_int_dat_o[5] ,
    \wbd_int_dat_o[4] ,
    \wbd_int_dat_o[3] ,
    \wbd_int_dat_o[2] ,
    \wbd_int_dat_o[1] ,
    \wbd_int_dat_o[0] }),
    .wbs_dat_o({\wbd_int_dat_i[31] ,
    \wbd_int_dat_i[30] ,
    \wbd_int_dat_i[29] ,
    \wbd_int_dat_i[28] ,
    \wbd_int_dat_i[27] ,
    \wbd_int_dat_i[26] ,
    \wbd_int_dat_i[25] ,
    \wbd_int_dat_i[24] ,
    \wbd_int_dat_i[23] ,
    \wbd_int_dat_i[22] ,
    \wbd_int_dat_i[21] ,
    \wbd_int_dat_i[20] ,
    \wbd_int_dat_i[19] ,
    \wbd_int_dat_i[18] ,
    \wbd_int_dat_i[17] ,
    \wbd_int_dat_i[16] ,
    \wbd_int_dat_i[15] ,
    \wbd_int_dat_i[14] ,
    \wbd_int_dat_i[13] ,
    \wbd_int_dat_i[12] ,
    \wbd_int_dat_i[11] ,
    \wbd_int_dat_i[10] ,
    \wbd_int_dat_i[9] ,
    \wbd_int_dat_i[8] ,
    \wbd_int_dat_i[7] ,
    \wbd_int_dat_i[6] ,
    \wbd_int_dat_i[5] ,
    \wbd_int_dat_i[4] ,
    \wbd_int_dat_i[3] ,
    \wbd_int_dat_i[2] ,
    \wbd_int_dat_i[1] ,
    \wbd_int_dat_i[0] }),
    .wbs_sel_o({\wbd_int_sel_i[3] ,
    \wbd_int_sel_i[2] ,
    \wbd_int_sel_i[1] ,
    \wbd_int_sel_i[0] }));
endmodule
